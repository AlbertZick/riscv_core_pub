module prim_ff_cl(
  input         clock,
  input         reset,
  output [19:0] io_q_op, 
  output [4:0]  io_q_dest, 
  output [4:0]  io_q_qj, 
  output [4:0]  io_q_qk, 
  output [31:0] io_q_a, 
  output [31:0] io_q_vj, 
  output [31:0] io_q_vk, 
  output        io_q_busy, 
  input  [19:0] io_d_op, 
  input  [4:0]  io_d_dest, 
  input  [4:0]  io_d_qj, 
  input  [4:0]  io_d_qk, 
  input  [31:0] io_d_a, 
  input  [31:0] io_d_vj, 
  input  [31:0] io_d_vk, 
  input         io_d_busy, 
  input         io_clear 
);
  reg [19:0] m_reg_op; 
  reg [4:0] m_reg_dest; 
  reg [4:0] m_reg_qj; 
  reg [4:0] m_reg_qk; 
  reg [31:0] m_reg_a; 
  reg [31:0] m_reg_vj; 
  reg [31:0] m_reg_vk; 
  reg  m_reg_busy; 
  assign io_q_op = m_reg_op; 
  assign io_q_dest = m_reg_dest; 
  assign io_q_qj = m_reg_qj; 
  assign io_q_qk = m_reg_qk; 
  assign io_q_a = m_reg_a; 
  assign io_q_vj = m_reg_vj; 
  assign io_q_vk = m_reg_vk; 
  assign io_q_busy = m_reg_busy; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_op <= 20'h0; 
    end else if (io_clear) begin 
      m_reg_op <= 20'h0;
    end else begin
      m_reg_op <= io_d_op;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_dest <= 5'h0; 
    end else if (io_clear) begin 
      m_reg_dest <= 5'h0;
    end else begin
      m_reg_dest <= io_d_dest;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_qj <= 5'h0; 
    end else if (io_clear) begin 
      m_reg_qj <= 5'h0;
    end else begin
      m_reg_qj <= io_d_qj;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_qk <= 5'h0; 
    end else if (io_clear) begin 
      m_reg_qk <= 5'h0;
    end else begin
      m_reg_qk <= io_d_qk;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_a <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_a <= 32'h0;
    end else begin
      m_reg_a <= io_d_a;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_vj <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_vj <= 32'h0;
    end else begin
      m_reg_vj <= io_d_vj;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_vk <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_vk <= 32'h0;
    end else begin
      m_reg_vk <= io_d_vk;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_busy <= 1'h0; 
    end else if (io_clear) begin 
      m_reg_busy <= 1'h0;
    end else begin
      m_reg_busy <= io_d_busy;
    end
  end
endmodule
module prim_ff_cl_4(
  input        clock,
  input        reset,
  output [3:0] io_q, 
  input  [3:0] io_d, 
  input        io_clear 
);
  reg [3:0] m_reg; 
  assign io_q = m_reg; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg <= 4'hf; 
    end else if (io_clear) begin 
      m_reg <= 4'hf;
    end else begin
      m_reg <= io_d;
    end
  end
endmodule
module integer_RS(
  input          clock,
  input          reset,
  input          io_clear, 
  input          io_enq, 
  input  [131:0] io_enq_data, 
  input          io_deq, 
  input  [3:0]   io_deq_cond, 
  output [131:0] io_deq_data, 
  output         io_empty, 
  output         io_full, 
  output [527:0] io_queue_data, 
  input  [3:0]   io_update_entry, 
  input  [527:0] io_update_entry_data 
);
  wire  FFs_0_clock; 
  wire  FFs_0_reset; 
  wire [19:0] FFs_0_io_q_op; 
  wire [4:0] FFs_0_io_q_dest; 
  wire [4:0] FFs_0_io_q_qj; 
  wire [4:0] FFs_0_io_q_qk; 
  wire [31:0] FFs_0_io_q_a; 
  wire [31:0] FFs_0_io_q_vj; 
  wire [31:0] FFs_0_io_q_vk; 
  wire  FFs_0_io_q_busy; 
  wire [19:0] FFs_0_io_d_op; 
  wire [4:0] FFs_0_io_d_dest; 
  wire [4:0] FFs_0_io_d_qj; 
  wire [4:0] FFs_0_io_d_qk; 
  wire [31:0] FFs_0_io_d_a; 
  wire [31:0] FFs_0_io_d_vj; 
  wire [31:0] FFs_0_io_d_vk; 
  wire  FFs_0_io_d_busy; 
  wire  FFs_0_io_clear; 
  wire  FFs_1_clock; 
  wire  FFs_1_reset; 
  wire [19:0] FFs_1_io_q_op; 
  wire [4:0] FFs_1_io_q_dest; 
  wire [4:0] FFs_1_io_q_qj; 
  wire [4:0] FFs_1_io_q_qk; 
  wire [31:0] FFs_1_io_q_a; 
  wire [31:0] FFs_1_io_q_vj; 
  wire [31:0] FFs_1_io_q_vk; 
  wire  FFs_1_io_q_busy; 
  wire [19:0] FFs_1_io_d_op; 
  wire [4:0] FFs_1_io_d_dest; 
  wire [4:0] FFs_1_io_d_qj; 
  wire [4:0] FFs_1_io_d_qk; 
  wire [31:0] FFs_1_io_d_a; 
  wire [31:0] FFs_1_io_d_vj; 
  wire [31:0] FFs_1_io_d_vk; 
  wire  FFs_1_io_d_busy; 
  wire  FFs_1_io_clear; 
  wire  FFs_2_clock; 
  wire  FFs_2_reset; 
  wire [19:0] FFs_2_io_q_op; 
  wire [4:0] FFs_2_io_q_dest; 
  wire [4:0] FFs_2_io_q_qj; 
  wire [4:0] FFs_2_io_q_qk; 
  wire [31:0] FFs_2_io_q_a; 
  wire [31:0] FFs_2_io_q_vj; 
  wire [31:0] FFs_2_io_q_vk; 
  wire  FFs_2_io_q_busy; 
  wire [19:0] FFs_2_io_d_op; 
  wire [4:0] FFs_2_io_d_dest; 
  wire [4:0] FFs_2_io_d_qj; 
  wire [4:0] FFs_2_io_d_qk; 
  wire [31:0] FFs_2_io_d_a; 
  wire [31:0] FFs_2_io_d_vj; 
  wire [31:0] FFs_2_io_d_vk; 
  wire  FFs_2_io_d_busy; 
  wire  FFs_2_io_clear; 
  wire  FFs_3_clock; 
  wire  FFs_3_reset; 
  wire [19:0] FFs_3_io_q_op; 
  wire [4:0] FFs_3_io_q_dest; 
  wire [4:0] FFs_3_io_q_qj; 
  wire [4:0] FFs_3_io_q_qk; 
  wire [31:0] FFs_3_io_q_a; 
  wire [31:0] FFs_3_io_q_vj; 
  wire [31:0] FFs_3_io_q_vk; 
  wire  FFs_3_io_q_busy; 
  wire [19:0] FFs_3_io_d_op; 
  wire [4:0] FFs_3_io_d_dest; 
  wire [4:0] FFs_3_io_d_qj; 
  wire [4:0] FFs_3_io_d_qk; 
  wire [31:0] FFs_3_io_d_a; 
  wire [31:0] FFs_3_io_d_vj; 
  wire [31:0] FFs_3_io_d_vk; 
  wire  FFs_3_io_d_busy; 
  wire  FFs_3_io_clear; 
  wire  mEntryEmpty_clock; 
  wire  mEntryEmpty_reset; 
  wire [3:0] mEntryEmpty_io_q; 
  wire [3:0] mEntryEmpty_io_d; 
  wire  mEntryEmpty_io_clear; 
  wire  _io_full_T = |mEntryEmpty_io_q; 
  wire [31:0] FFs_io_0_q_vk = FFs_0_io_q_vk; 
  wire  FFs_io_0_q_busy = FFs_0_io_q_busy; 
  wire [31:0] FFs_io_0_q_a = FFs_0_io_q_a; 
  wire [31:0] FFs_io_0_q_vj = FFs_0_io_q_vj; 
  wire [4:0] FFs_io_0_q_qj = FFs_0_io_q_qj; 
  wire [4:0] FFs_io_0_q_qk = FFs_0_io_q_qk; 
  wire [19:0] FFs_io_0_q_op = FFs_0_io_q_op; 
  wire [4:0] FFs_io_0_q_dest = FFs_0_io_q_dest; 
  wire [131:0] io_queue_data_lo_lo = {FFs_io_0_q_op,FFs_io_0_q_dest,FFs_io_0_q_qj,FFs_io_0_q_qk,FFs_io_0_q_a,
    FFs_io_0_q_vj,FFs_io_0_q_vk,FFs_io_0_q_busy}; 
  wire [31:0] FFs_io_1_q_vk = FFs_1_io_q_vk; 
  wire  FFs_io_1_q_busy = FFs_1_io_q_busy; 
  wire [31:0] FFs_io_1_q_a = FFs_1_io_q_a; 
  wire [31:0] FFs_io_1_q_vj = FFs_1_io_q_vj; 
  wire [4:0] FFs_io_1_q_qj = FFs_1_io_q_qj; 
  wire [4:0] FFs_io_1_q_qk = FFs_1_io_q_qk; 
  wire [19:0] FFs_io_1_q_op = FFs_1_io_q_op; 
  wire [4:0] FFs_io_1_q_dest = FFs_1_io_q_dest; 
  wire [263:0] io_queue_data_lo = {FFs_io_1_q_op,FFs_io_1_q_dest,FFs_io_1_q_qj,FFs_io_1_q_qk,FFs_io_1_q_a,FFs_io_1_q_vj,
    FFs_io_1_q_vk,FFs_io_1_q_busy,io_queue_data_lo_lo}; 
  wire [31:0] FFs_io_2_q_vk = FFs_2_io_q_vk; 
  wire  FFs_io_2_q_busy = FFs_2_io_q_busy; 
  wire [31:0] FFs_io_2_q_a = FFs_2_io_q_a; 
  wire [31:0] FFs_io_2_q_vj = FFs_2_io_q_vj; 
  wire [4:0] FFs_io_2_q_qj = FFs_2_io_q_qj; 
  wire [4:0] FFs_io_2_q_qk = FFs_2_io_q_qk; 
  wire [19:0] FFs_io_2_q_op = FFs_2_io_q_op; 
  wire [4:0] FFs_io_2_q_dest = FFs_2_io_q_dest; 
  wire [131:0] io_queue_data_hi_lo = {FFs_io_2_q_op,FFs_io_2_q_dest,FFs_io_2_q_qj,FFs_io_2_q_qk,FFs_io_2_q_a,
    FFs_io_2_q_vj,FFs_io_2_q_vk,FFs_io_2_q_busy}; 
  wire [31:0] FFs_io_3_q_vk = FFs_3_io_q_vk; 
  wire  FFs_io_3_q_busy = FFs_3_io_q_busy; 
  wire [31:0] FFs_io_3_q_a = FFs_3_io_q_a; 
  wire [31:0] FFs_io_3_q_vj = FFs_3_io_q_vj; 
  wire [4:0] FFs_io_3_q_qj = FFs_3_io_q_qj; 
  wire [4:0] FFs_io_3_q_qk = FFs_3_io_q_qk; 
  wire [19:0] FFs_io_3_q_op = FFs_3_io_q_op; 
  wire [4:0] FFs_io_3_q_dest = FFs_3_io_q_dest; 
  wire [263:0] io_queue_data_hi = {FFs_io_3_q_op,FFs_io_3_q_dest,FFs_io_3_q_qj,FFs_io_3_q_qk,FFs_io_3_q_a,FFs_io_3_q_vj,
    FFs_io_3_q_vk,FFs_io_3_q_busy,io_queue_data_hi_lo}; 
  wire  _oneHotDeqCond_0_T_1 = ~mEntryEmpty_io_q[0]; 
  wire  oneHotDeqCond_0 = io_deq & ~mEntryEmpty_io_q[0] & io_deq_cond[0]; 
  wire  oneHotEnq_0 = io_enq & mEntryEmpty_io_q[0]; 
  wire  updateEntryVl_0 = io_update_entry[0] & _oneHotDeqCond_0_T_1; 
  wire  _GEN_0 = oneHotEnq_0 ? io_enq_data[0] : FFs_io_0_q_busy; 
  wire [31:0] _GEN_1 = oneHotEnq_0 ? io_enq_data[32:1] : FFs_io_0_q_vk; 
  wire [31:0] _GEN_2 = oneHotEnq_0 ? io_enq_data[64:33] : FFs_io_0_q_vj; 
  wire [31:0] _GEN_3 = oneHotEnq_0 ? io_enq_data[96:65] : FFs_io_0_q_a; 
  wire [4:0] _GEN_4 = oneHotEnq_0 ? io_enq_data[101:97] : FFs_io_0_q_qk; 
  wire [4:0] _GEN_5 = oneHotEnq_0 ? io_enq_data[106:102] : FFs_io_0_q_qj; 
  wire [4:0] _GEN_6 = oneHotEnq_0 ? io_enq_data[111:107] : FFs_io_0_q_dest; 
  wire [19:0] _GEN_7 = oneHotEnq_0 ? io_enq_data[131:112] : FFs_io_0_q_op; 
  wire  updatedData_0_busy = updateEntryVl_0 ? io_update_entry_data[0] : _GEN_0; 
  wire [31:0] updatedData_0_vk = updateEntryVl_0 ? io_update_entry_data[32:1] : _GEN_1; 
  wire [31:0] updatedData_0_vj = updateEntryVl_0 ? io_update_entry_data[64:33] : _GEN_2; 
  wire [31:0] updatedData_0_a = updateEntryVl_0 ? io_update_entry_data[96:65] : _GEN_3; 
  wire [4:0] updatedData_0_qk = updateEntryVl_0 ? io_update_entry_data[101:97] : _GEN_4; 
  wire [4:0] updatedData_0_qj = updateEntryVl_0 ? io_update_entry_data[106:102] : _GEN_5; 
  wire [4:0] updatedData_0_dest = updateEntryVl_0 ? io_update_entry_data[111:107] : _GEN_6; 
  wire [19:0] updatedData_0_op = updateEntryVl_0 ? io_update_entry_data[131:112] : _GEN_7; 
  wire  _oneHotDeqCond_1_T_1 = ~mEntryEmpty_io_q[1]; 
  wire  _oneHotDeqCond_1_T_7 = ~(|io_deq_cond[0]); 
  wire  oneHotDeqCond_1 = io_deq & ~mEntryEmpty_io_q[1] & io_deq_cond[1] & _oneHotDeqCond_1_T_7; 
  wire  oneHotEnq_1 = io_enq & mEntryEmpty_io_q[1] & ~(|mEntryEmpty_io_q[0]); 
  wire  updateEntryVl_1 = io_update_entry[1] & _oneHotDeqCond_1_T_1; 
  wire  _GEN_16 = oneHotEnq_1 ? io_enq_data[0] : FFs_io_1_q_busy; 
  wire [31:0] _GEN_17 = oneHotEnq_1 ? io_enq_data[32:1] : FFs_io_1_q_vk; 
  wire [31:0] _GEN_18 = oneHotEnq_1 ? io_enq_data[64:33] : FFs_io_1_q_vj; 
  wire [31:0] _GEN_19 = oneHotEnq_1 ? io_enq_data[96:65] : FFs_io_1_q_a; 
  wire [4:0] _GEN_20 = oneHotEnq_1 ? io_enq_data[101:97] : FFs_io_1_q_qk; 
  wire [4:0] _GEN_21 = oneHotEnq_1 ? io_enq_data[106:102] : FFs_io_1_q_qj; 
  wire [4:0] _GEN_22 = oneHotEnq_1 ? io_enq_data[111:107] : FFs_io_1_q_dest; 
  wire [19:0] _GEN_23 = oneHotEnq_1 ? io_enq_data[131:112] : FFs_io_1_q_op; 
  wire  updatedData_1_busy = updateEntryVl_1 ? io_update_entry_data[132] : _GEN_16; 
  wire [31:0] updatedData_1_vk = updateEntryVl_1 ? io_update_entry_data[164:133] : _GEN_17; 
  wire [31:0] updatedData_1_vj = updateEntryVl_1 ? io_update_entry_data[196:165] : _GEN_18; 
  wire [31:0] updatedData_1_a = updateEntryVl_1 ? io_update_entry_data[228:197] : _GEN_19; 
  wire [4:0] updatedData_1_qk = updateEntryVl_1 ? io_update_entry_data[233:229] : _GEN_20; 
  wire [4:0] updatedData_1_qj = updateEntryVl_1 ? io_update_entry_data[238:234] : _GEN_21; 
  wire [4:0] updatedData_1_dest = updateEntryVl_1 ? io_update_entry_data[243:239] : _GEN_22; 
  wire [19:0] updatedData_1_op = updateEntryVl_1 ? io_update_entry_data[263:244] : _GEN_23; 
  wire  _oneHotDeqCond_2_T_1 = ~mEntryEmpty_io_q[2]; 
  wire  _oneHotDeqCond_2_T_7 = ~(|io_deq_cond[1:0]); 
  wire  oneHotDeqCond_2 = io_deq & ~mEntryEmpty_io_q[2] & io_deq_cond[2] & _oneHotDeqCond_2_T_7; 
  wire  oneHotEnq_2 = io_enq & mEntryEmpty_io_q[2] & ~(|mEntryEmpty_io_q[1:0]); 
  wire  updateEntryVl_2 = io_update_entry[2] & _oneHotDeqCond_2_T_1; 
  wire  _GEN_32 = oneHotEnq_2 ? io_enq_data[0] : FFs_io_2_q_busy; 
  wire [31:0] _GEN_33 = oneHotEnq_2 ? io_enq_data[32:1] : FFs_io_2_q_vk; 
  wire [31:0] _GEN_34 = oneHotEnq_2 ? io_enq_data[64:33] : FFs_io_2_q_vj; 
  wire [31:0] _GEN_35 = oneHotEnq_2 ? io_enq_data[96:65] : FFs_io_2_q_a; 
  wire [4:0] _GEN_36 = oneHotEnq_2 ? io_enq_data[101:97] : FFs_io_2_q_qk; 
  wire [4:0] _GEN_37 = oneHotEnq_2 ? io_enq_data[106:102] : FFs_io_2_q_qj; 
  wire [4:0] _GEN_38 = oneHotEnq_2 ? io_enq_data[111:107] : FFs_io_2_q_dest; 
  wire [19:0] _GEN_39 = oneHotEnq_2 ? io_enq_data[131:112] : FFs_io_2_q_op; 
  wire  updatedData_2_busy = updateEntryVl_2 ? io_update_entry_data[264] : _GEN_32; 
  wire [31:0] updatedData_2_vk = updateEntryVl_2 ? io_update_entry_data[296:265] : _GEN_33; 
  wire [31:0] updatedData_2_vj = updateEntryVl_2 ? io_update_entry_data[328:297] : _GEN_34; 
  wire [31:0] updatedData_2_a = updateEntryVl_2 ? io_update_entry_data[360:329] : _GEN_35; 
  wire [4:0] updatedData_2_qk = updateEntryVl_2 ? io_update_entry_data[365:361] : _GEN_36; 
  wire [4:0] updatedData_2_qj = updateEntryVl_2 ? io_update_entry_data[370:366] : _GEN_37; 
  wire [4:0] updatedData_2_dest = updateEntryVl_2 ? io_update_entry_data[375:371] : _GEN_38; 
  wire [19:0] updatedData_2_op = updateEntryVl_2 ? io_update_entry_data[395:376] : _GEN_39; 
  wire  _oneHotDeqCond_3_T_1 = ~mEntryEmpty_io_q[3]; 
  wire  _oneHotDeqCond_3_T_7 = ~(|io_deq_cond[2:0]); 
  wire  oneHotDeqCond_3 = io_deq & ~mEntryEmpty_io_q[3] & io_deq_cond[3] & _oneHotDeqCond_3_T_7; 
  wire  oneHotEnq_3 = io_enq & mEntryEmpty_io_q[3] & ~(|mEntryEmpty_io_q[2:0]); 
  wire  updateEntryVl_3 = io_update_entry[3] & _oneHotDeqCond_3_T_1; 
  wire  _GEN_48 = oneHotEnq_3 ? io_enq_data[0] : FFs_io_3_q_busy; 
  wire [31:0] _GEN_49 = oneHotEnq_3 ? io_enq_data[32:1] : FFs_io_3_q_vk; 
  wire [31:0] _GEN_50 = oneHotEnq_3 ? io_enq_data[64:33] : FFs_io_3_q_vj; 
  wire [31:0] _GEN_51 = oneHotEnq_3 ? io_enq_data[96:65] : FFs_io_3_q_a; 
  wire [4:0] _GEN_52 = oneHotEnq_3 ? io_enq_data[101:97] : FFs_io_3_q_qk; 
  wire [4:0] _GEN_53 = oneHotEnq_3 ? io_enq_data[106:102] : FFs_io_3_q_qj; 
  wire [4:0] _GEN_54 = oneHotEnq_3 ? io_enq_data[111:107] : FFs_io_3_q_dest; 
  wire [19:0] _GEN_55 = oneHotEnq_3 ? io_enq_data[131:112] : FFs_io_3_q_op; 
  wire  updatedData_3_busy = updateEntryVl_3 ? io_update_entry_data[396] : _GEN_48; 
  wire [31:0] updatedData_3_vk = updateEntryVl_3 ? io_update_entry_data[428:397] : _GEN_49; 
  wire [31:0] updatedData_3_vj = updateEntryVl_3 ? io_update_entry_data[460:429] : _GEN_50; 
  wire [31:0] updatedData_3_a = updateEntryVl_3 ? io_update_entry_data[492:461] : _GEN_51; 
  wire [4:0] updatedData_3_qk = updateEntryVl_3 ? io_update_entry_data[497:493] : _GEN_52; 
  wire [4:0] updatedData_3_qj = updateEntryVl_3 ? io_update_entry_data[502:498] : _GEN_53; 
  wire [4:0] updatedData_3_dest = updateEntryVl_3 ? io_update_entry_data[507:503] : _GEN_54; 
  wire [19:0] updatedData_3_op = updateEntryVl_3 ? io_update_entry_data[527:508] : _GEN_55; 
  wire [1:0] _GEN_66 = oneHotDeqCond_2 ? 2'h2 : {{1'd0}, oneHotDeqCond_1}; 
  wire [1:0] oneHotDeqCond_idx = oneHotDeqCond_3 ? 2'h3 : _GEN_66; 
  wire  enqVl = io_enq & _io_full_T; 
  wire [31:0] _GEN_69 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_vk : FFs_io_0_q_vk; 
  wire [31:0] _GEN_70 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_vk : _GEN_69; 
  wire [31:0] _GEN_71 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_vk : _GEN_70; 
  wire  _GEN_73 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_busy : FFs_io_0_q_busy; 
  wire  _GEN_74 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_busy : _GEN_73; 
  wire  _GEN_75 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_busy : _GEN_74; 
  wire [31:0] _GEN_77 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_a : FFs_io_0_q_a; 
  wire [31:0] _GEN_78 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_a : _GEN_77; 
  wire [31:0] _GEN_79 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_a : _GEN_78; 
  wire [31:0] _GEN_81 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_vj : FFs_io_0_q_vj; 
  wire [31:0] _GEN_82 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_vj : _GEN_81; 
  wire [31:0] _GEN_83 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_vj : _GEN_82; 
  wire [4:0] _GEN_85 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_qj : FFs_io_0_q_qj; 
  wire [4:0] _GEN_86 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_qj : _GEN_85; 
  wire [4:0] _GEN_87 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_qj : _GEN_86; 
  wire [4:0] _GEN_89 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_qk : FFs_io_0_q_qk; 
  wire [4:0] _GEN_90 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_qk : _GEN_89; 
  wire [4:0] _GEN_91 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_qk : _GEN_90; 
  wire [19:0] _GEN_93 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_op : FFs_io_0_q_op; 
  wire [19:0] _GEN_94 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_op : _GEN_93; 
  wire [19:0] _GEN_95 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_op : _GEN_94; 
  wire [4:0] _GEN_97 = 2'h1 == oneHotDeqCond_idx ? FFs_io_1_q_dest : FFs_io_0_q_dest; 
  wire [4:0] _GEN_98 = 2'h2 == oneHotDeqCond_idx ? FFs_io_2_q_dest : _GEN_97; 
  wire [4:0] _GEN_99 = 2'h3 == oneHotDeqCond_idx ? FFs_io_3_q_dest : _GEN_98; 
  wire [131:0] _io_deq_data_T = {_GEN_95,_GEN_99,_GEN_87,_GEN_91,_GEN_79,_GEN_83,_GEN_71,_GEN_75}; 
  wire [3:0] _T_16 = {oneHotDeqCond_3,oneHotDeqCond_2,oneHotDeqCond_1,oneHotDeqCond_0}; 
  wire  _T_20 = ~enqVl; 
  wire [3:0] _mEntryEmpty_io_d_T_1 = {1'h1,mEntryEmpty_io_q[3:1]}; 
  wire [3:0] _GEN_100 = ~enqVl ? _mEntryEmpty_io_d_T_1 : mEntryEmpty_io_q; 
  wire  _GEN_101 = &mEntryEmpty_io_q[3:1] & _T_20 | io_clear; 
  wire  _GEN_102 = 2'h0 == oneHotDeqCond_idx ? _GEN_101 : io_clear; 
  wire  _GEN_111 = 2'h0 < oneHotDeqCond_idx ? io_clear : _GEN_102; 
  wire  _GEN_112 = &mEntryEmpty_io_q[3:2] & _T_20 | io_clear; 
  wire  _GEN_113 = 2'h1 == oneHotDeqCond_idx ? _GEN_112 : io_clear; 
  wire  _GEN_114 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_busy : updatedData_1_busy; 
  wire [31:0] _GEN_115 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_vk : updatedData_1_vk; 
  wire [31:0] _GEN_116 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_vj : updatedData_1_vj; 
  wire [31:0] _GEN_117 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_a : updatedData_1_a; 
  wire [4:0] _GEN_118 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_qk : updatedData_1_qk; 
  wire [4:0] _GEN_119 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_qj : updatedData_1_qj; 
  wire [4:0] _GEN_120 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_dest : updatedData_1_dest; 
  wire [19:0] _GEN_121 = 2'h1 == oneHotDeqCond_idx ? updatedData_0_op : updatedData_1_op; 
  wire  _GEN_130 = 2'h1 < oneHotDeqCond_idx ? io_clear : _GEN_113; 
  wire  _GEN_131 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_busy : _GEN_114; 
  wire [31:0] _GEN_132 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_vk : _GEN_115; 
  wire [31:0] _GEN_133 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_vj : _GEN_116; 
  wire [31:0] _GEN_134 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_a : _GEN_117; 
  wire [4:0] _GEN_135 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_qk : _GEN_118; 
  wire [4:0] _GEN_136 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_qj : _GEN_119; 
  wire [4:0] _GEN_137 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_dest : _GEN_120; 
  wire [19:0] _GEN_138 = 2'h1 < oneHotDeqCond_idx ? updatedData_0_op : _GEN_121; 
  wire  _GEN_139 = &mEntryEmpty_io_q[3] & _T_20 | io_clear; 
  wire  _GEN_140 = 2'h2 == oneHotDeqCond_idx ? _GEN_139 : io_clear; 
  wire  _GEN_141 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_busy : updatedData_2_busy; 
  wire [31:0] _GEN_142 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_vk : updatedData_2_vk; 
  wire [31:0] _GEN_143 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_vj : updatedData_2_vj; 
  wire [31:0] _GEN_144 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_a : updatedData_2_a; 
  wire [4:0] _GEN_145 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_qk : updatedData_2_qk; 
  wire [4:0] _GEN_146 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_qj : updatedData_2_qj; 
  wire [4:0] _GEN_147 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_dest : updatedData_2_dest; 
  wire [19:0] _GEN_148 = 2'h2 == oneHotDeqCond_idx ? updatedData_1_op : updatedData_2_op; 
  wire  _GEN_157 = 2'h2 < oneHotDeqCond_idx ? io_clear : _GEN_140; 
  wire  _GEN_158 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_busy : _GEN_141; 
  wire [31:0] _GEN_159 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_vk : _GEN_142; 
  wire [31:0] _GEN_160 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_vj : _GEN_143; 
  wire [31:0] _GEN_161 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_a : _GEN_144; 
  wire [4:0] _GEN_162 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_qk : _GEN_145; 
  wire [4:0] _GEN_163 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_qj : _GEN_146; 
  wire [4:0] _GEN_164 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_dest : _GEN_147; 
  wire [19:0] _GEN_165 = 2'h2 < oneHotDeqCond_idx ? updatedData_1_op : _GEN_148; 
  wire  _GEN_166 = _T_20 | io_clear; 
  wire  _GEN_167 = 2'h3 == oneHotDeqCond_idx | _GEN_166; 
  wire  _GEN_168 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_busy : updatedData_3_busy; 
  wire [31:0] _GEN_169 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_vk : updatedData_3_vk; 
  wire [31:0] _GEN_170 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_vj : updatedData_3_vj; 
  wire [31:0] _GEN_171 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_a : updatedData_3_a; 
  wire [4:0] _GEN_172 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_qk : updatedData_3_qk; 
  wire [4:0] _GEN_173 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_qj : updatedData_3_qj; 
  wire [4:0] _GEN_174 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_dest : updatedData_3_dest; 
  wire [19:0] _GEN_175 = 2'h3 == oneHotDeqCond_idx ? updatedData_2_op : updatedData_3_op; 
  wire [3:0] _mEntryEmpty_io_d_T_3 = {mEntryEmpty_io_q[3:1],1'h0}; 
  wire [3:0] _GEN_193 = oneHotEnq_0 ? _mEntryEmpty_io_d_T_3 : mEntryEmpty_io_q; 
  wire [3:0] _GEN_194 = updateEntryVl_0 ? mEntryEmpty_io_q : _GEN_193; 
  wire [3:0] _mEntryEmpty_io_d_T_6 = {mEntryEmpty_io_q[3:2],1'h0,mEntryEmpty_io_q[0]}; 
  wire [3:0] _GEN_195 = oneHotEnq_1 ? _mEntryEmpty_io_d_T_6 : _GEN_194; 
  wire [3:0] _GEN_196 = updateEntryVl_1 ? _GEN_194 : _GEN_195; 
  wire [3:0] _mEntryEmpty_io_d_T_9 = {mEntryEmpty_io_q[3],1'h0,mEntryEmpty_io_q[1:0]}; 
  wire [3:0] _GEN_197 = oneHotEnq_2 ? _mEntryEmpty_io_d_T_9 : _GEN_196; 
  wire [3:0] _GEN_198 = updateEntryVl_2 ? _GEN_196 : _GEN_197; 
  wire [3:0] _mEntryEmpty_io_d_T_11 = {1'h0,mEntryEmpty_io_q[2:0]}; 
  wire [3:0] _GEN_199 = oneHotEnq_3 ? _mEntryEmpty_io_d_T_11 : _GEN_198; 
  wire [3:0] _GEN_200 = updateEntryVl_3 ? _GEN_198 : _GEN_199; 
  prim_ff_cl FFs_0 ( 
    .clock(FFs_0_clock),
    .reset(FFs_0_reset),
    .io_q_op(FFs_0_io_q_op),
    .io_q_dest(FFs_0_io_q_dest),
    .io_q_qj(FFs_0_io_q_qj),
    .io_q_qk(FFs_0_io_q_qk),
    .io_q_a(FFs_0_io_q_a),
    .io_q_vj(FFs_0_io_q_vj),
    .io_q_vk(FFs_0_io_q_vk),
    .io_q_busy(FFs_0_io_q_busy),
    .io_d_op(FFs_0_io_d_op),
    .io_d_dest(FFs_0_io_d_dest),
    .io_d_qj(FFs_0_io_d_qj),
    .io_d_qk(FFs_0_io_d_qk),
    .io_d_a(FFs_0_io_d_a),
    .io_d_vj(FFs_0_io_d_vj),
    .io_d_vk(FFs_0_io_d_vk),
    .io_d_busy(FFs_0_io_d_busy),
    .io_clear(FFs_0_io_clear)
  );
  prim_ff_cl FFs_1 ( 
    .clock(FFs_1_clock),
    .reset(FFs_1_reset),
    .io_q_op(FFs_1_io_q_op),
    .io_q_dest(FFs_1_io_q_dest),
    .io_q_qj(FFs_1_io_q_qj),
    .io_q_qk(FFs_1_io_q_qk),
    .io_q_a(FFs_1_io_q_a),
    .io_q_vj(FFs_1_io_q_vj),
    .io_q_vk(FFs_1_io_q_vk),
    .io_q_busy(FFs_1_io_q_busy),
    .io_d_op(FFs_1_io_d_op),
    .io_d_dest(FFs_1_io_d_dest),
    .io_d_qj(FFs_1_io_d_qj),
    .io_d_qk(FFs_1_io_d_qk),
    .io_d_a(FFs_1_io_d_a),
    .io_d_vj(FFs_1_io_d_vj),
    .io_d_vk(FFs_1_io_d_vk),
    .io_d_busy(FFs_1_io_d_busy),
    .io_clear(FFs_1_io_clear)
  );
  prim_ff_cl FFs_2 ( 
    .clock(FFs_2_clock),
    .reset(FFs_2_reset),
    .io_q_op(FFs_2_io_q_op),
    .io_q_dest(FFs_2_io_q_dest),
    .io_q_qj(FFs_2_io_q_qj),
    .io_q_qk(FFs_2_io_q_qk),
    .io_q_a(FFs_2_io_q_a),
    .io_q_vj(FFs_2_io_q_vj),
    .io_q_vk(FFs_2_io_q_vk),
    .io_q_busy(FFs_2_io_q_busy),
    .io_d_op(FFs_2_io_d_op),
    .io_d_dest(FFs_2_io_d_dest),
    .io_d_qj(FFs_2_io_d_qj),
    .io_d_qk(FFs_2_io_d_qk),
    .io_d_a(FFs_2_io_d_a),
    .io_d_vj(FFs_2_io_d_vj),
    .io_d_vk(FFs_2_io_d_vk),
    .io_d_busy(FFs_2_io_d_busy),
    .io_clear(FFs_2_io_clear)
  );
  prim_ff_cl FFs_3 ( 
    .clock(FFs_3_clock),
    .reset(FFs_3_reset),
    .io_q_op(FFs_3_io_q_op),
    .io_q_dest(FFs_3_io_q_dest),
    .io_q_qj(FFs_3_io_q_qj),
    .io_q_qk(FFs_3_io_q_qk),
    .io_q_a(FFs_3_io_q_a),
    .io_q_vj(FFs_3_io_q_vj),
    .io_q_vk(FFs_3_io_q_vk),
    .io_q_busy(FFs_3_io_q_busy),
    .io_d_op(FFs_3_io_d_op),
    .io_d_dest(FFs_3_io_d_dest),
    .io_d_qj(FFs_3_io_d_qj),
    .io_d_qk(FFs_3_io_d_qk),
    .io_d_a(FFs_3_io_d_a),
    .io_d_vj(FFs_3_io_d_vj),
    .io_d_vk(FFs_3_io_d_vk),
    .io_d_busy(FFs_3_io_d_busy),
    .io_clear(FFs_3_io_clear)
  );
  prim_ff_cl_4 mEntryEmpty ( 
    .clock(mEntryEmpty_clock),
    .reset(mEntryEmpty_reset),
    .io_q(mEntryEmpty_io_q),
    .io_d(mEntryEmpty_io_d),
    .io_clear(mEntryEmpty_io_clear)
  );
  assign io_deq_data = |_T_16 ? _io_deq_data_T : io_queue_data_lo_lo; 
  assign io_empty = &mEntryEmpty_io_q; 
  assign io_full = ~(|mEntryEmpty_io_q); 
  assign io_queue_data = {io_queue_data_hi,io_queue_data_lo}; 
  assign FFs_0_clock = clock;
  assign FFs_0_reset = reset;
  assign FFs_0_io_d_op = |_T_16 ? _GEN_138 : updatedData_0_op; 
  assign FFs_0_io_d_dest = |_T_16 ? _GEN_137 : updatedData_0_dest; 
  assign FFs_0_io_d_qj = |_T_16 ? _GEN_136 : updatedData_0_qj; 
  assign FFs_0_io_d_qk = |_T_16 ? _GEN_135 : updatedData_0_qk; 
  assign FFs_0_io_d_a = |_T_16 ? _GEN_134 : updatedData_0_a; 
  assign FFs_0_io_d_vj = |_T_16 ? _GEN_133 : updatedData_0_vj; 
  assign FFs_0_io_d_vk = |_T_16 ? _GEN_132 : updatedData_0_vk; 
  assign FFs_0_io_d_busy = |_T_16 ? _GEN_131 : updatedData_0_busy; 
  assign FFs_0_io_clear = |_T_16 ? _GEN_111 : io_clear; 
  assign FFs_1_clock = clock;
  assign FFs_1_reset = reset;
  assign FFs_1_io_d_op = |_T_16 ? _GEN_165 : updatedData_1_op; 
  assign FFs_1_io_d_dest = |_T_16 ? _GEN_164 : updatedData_1_dest; 
  assign FFs_1_io_d_qj = |_T_16 ? _GEN_163 : updatedData_1_qj; 
  assign FFs_1_io_d_qk = |_T_16 ? _GEN_162 : updatedData_1_qk; 
  assign FFs_1_io_d_a = |_T_16 ? _GEN_161 : updatedData_1_a; 
  assign FFs_1_io_d_vj = |_T_16 ? _GEN_160 : updatedData_1_vj; 
  assign FFs_1_io_d_vk = |_T_16 ? _GEN_159 : updatedData_1_vk; 
  assign FFs_1_io_d_busy = |_T_16 ? _GEN_158 : updatedData_1_busy; 
  assign FFs_1_io_clear = |_T_16 ? _GEN_130 : io_clear; 
  assign FFs_2_clock = clock;
  assign FFs_2_reset = reset;
  assign FFs_2_io_d_op = |_T_16 ? _GEN_175 : updatedData_2_op; 
  assign FFs_2_io_d_dest = |_T_16 ? _GEN_174 : updatedData_2_dest; 
  assign FFs_2_io_d_qj = |_T_16 ? _GEN_173 : updatedData_2_qj; 
  assign FFs_2_io_d_qk = |_T_16 ? _GEN_172 : updatedData_2_qk; 
  assign FFs_2_io_d_a = |_T_16 ? _GEN_171 : updatedData_2_a; 
  assign FFs_2_io_d_vj = |_T_16 ? _GEN_170 : updatedData_2_vj; 
  assign FFs_2_io_d_vk = |_T_16 ? _GEN_169 : updatedData_2_vk; 
  assign FFs_2_io_d_busy = |_T_16 ? _GEN_168 : updatedData_2_busy; 
  assign FFs_2_io_clear = |_T_16 ? _GEN_157 : io_clear; 
  assign FFs_3_clock = clock;
  assign FFs_3_reset = reset;
  assign FFs_3_io_d_op = updateEntryVl_3 ? io_update_entry_data[527:508] : _GEN_55; 
  assign FFs_3_io_d_dest = updateEntryVl_3 ? io_update_entry_data[507:503] : _GEN_54; 
  assign FFs_3_io_d_qj = updateEntryVl_3 ? io_update_entry_data[502:498] : _GEN_53; 
  assign FFs_3_io_d_qk = updateEntryVl_3 ? io_update_entry_data[497:493] : _GEN_52; 
  assign FFs_3_io_d_a = updateEntryVl_3 ? io_update_entry_data[492:461] : _GEN_51; 
  assign FFs_3_io_d_vj = updateEntryVl_3 ? io_update_entry_data[460:429] : _GEN_50; 
  assign FFs_3_io_d_vk = updateEntryVl_3 ? io_update_entry_data[428:397] : _GEN_49; 
  assign FFs_3_io_d_busy = updateEntryVl_3 ? io_update_entry_data[396] : _GEN_48; 
  assign FFs_3_io_clear = |_T_16 ? _GEN_167 : io_clear; 
  assign mEntryEmpty_clock = clock;
  assign mEntryEmpty_reset = reset;
  assign mEntryEmpty_io_d = |_T_16 ? _GEN_100 : _GEN_200; 
  assign mEntryEmpty_io_clear = io_clear; 
endmodule
module prim_ff_cl_5(
  input        clock,
  input        reset,
  output [1:0] io_q, 
  input  [1:0] io_d, 
  input        io_clear 
);
  reg [1:0] m_reg; 
  assign io_q = m_reg; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg <= 2'h0; 
    end else if (io_clear) begin 
      m_reg <= 2'h0;
    end else begin
      m_reg <= io_d;
    end
  end
endmodule
module FIFO(
  input          clock,
  input          reset,
  input          io_clear, 
  input          io_enq, 
  input  [131:0] io_enq_data, 
  output [1:0]   io_enq_idx, 
  input          io_deq, 
  output [131:0] io_deq_data, 
  output [1:0]   io_deq_idx, 
  output         io_empty, 
  output         io_full, 
  output [527:0] io_queue_data, 
  input  [3:0]   io_update_entry, 
  input  [527:0] io_update_entry_data 
);
  wire  h_ptr_clock; 
  wire  h_ptr_reset; 
  wire [1:0] h_ptr_io_q; 
  wire [1:0] h_ptr_io_d; 
  wire  h_ptr_io_clear; 
  wire  t_ptr_clock; 
  wire  t_ptr_reset; 
  wire [1:0] t_ptr_io_q; 
  wire [1:0] t_ptr_io_d; 
  wire  t_ptr_io_clear; 
  wire  FFs_0_clock; 
  wire  FFs_0_reset; 
  wire [19:0] FFs_0_io_q_op; 
  wire [4:0] FFs_0_io_q_dest; 
  wire [4:0] FFs_0_io_q_qj; 
  wire [4:0] FFs_0_io_q_qk; 
  wire [31:0] FFs_0_io_q_a; 
  wire [31:0] FFs_0_io_q_vj; 
  wire [31:0] FFs_0_io_q_vk; 
  wire  FFs_0_io_q_busy; 
  wire [19:0] FFs_0_io_d_op; 
  wire [4:0] FFs_0_io_d_dest; 
  wire [4:0] FFs_0_io_d_qj; 
  wire [4:0] FFs_0_io_d_qk; 
  wire [31:0] FFs_0_io_d_a; 
  wire [31:0] FFs_0_io_d_vj; 
  wire [31:0] FFs_0_io_d_vk; 
  wire  FFs_0_io_d_busy; 
  wire  FFs_0_io_clear; 
  wire  FFs_1_clock; 
  wire  FFs_1_reset; 
  wire [19:0] FFs_1_io_q_op; 
  wire [4:0] FFs_1_io_q_dest; 
  wire [4:0] FFs_1_io_q_qj; 
  wire [4:0] FFs_1_io_q_qk; 
  wire [31:0] FFs_1_io_q_a; 
  wire [31:0] FFs_1_io_q_vj; 
  wire [31:0] FFs_1_io_q_vk; 
  wire  FFs_1_io_q_busy; 
  wire [19:0] FFs_1_io_d_op; 
  wire [4:0] FFs_1_io_d_dest; 
  wire [4:0] FFs_1_io_d_qj; 
  wire [4:0] FFs_1_io_d_qk; 
  wire [31:0] FFs_1_io_d_a; 
  wire [31:0] FFs_1_io_d_vj; 
  wire [31:0] FFs_1_io_d_vk; 
  wire  FFs_1_io_d_busy; 
  wire  FFs_1_io_clear; 
  wire  FFs_2_clock; 
  wire  FFs_2_reset; 
  wire [19:0] FFs_2_io_q_op; 
  wire [4:0] FFs_2_io_q_dest; 
  wire [4:0] FFs_2_io_q_qj; 
  wire [4:0] FFs_2_io_q_qk; 
  wire [31:0] FFs_2_io_q_a; 
  wire [31:0] FFs_2_io_q_vj; 
  wire [31:0] FFs_2_io_q_vk; 
  wire  FFs_2_io_q_busy; 
  wire [19:0] FFs_2_io_d_op; 
  wire [4:0] FFs_2_io_d_dest; 
  wire [4:0] FFs_2_io_d_qj; 
  wire [4:0] FFs_2_io_d_qk; 
  wire [31:0] FFs_2_io_d_a; 
  wire [31:0] FFs_2_io_d_vj; 
  wire [31:0] FFs_2_io_d_vk; 
  wire  FFs_2_io_d_busy; 
  wire  FFs_2_io_clear; 
  wire  FFs_3_clock; 
  wire  FFs_3_reset; 
  wire [19:0] FFs_3_io_q_op; 
  wire [4:0] FFs_3_io_q_dest; 
  wire [4:0] FFs_3_io_q_qj; 
  wire [4:0] FFs_3_io_q_qk; 
  wire [31:0] FFs_3_io_q_a; 
  wire [31:0] FFs_3_io_q_vj; 
  wire [31:0] FFs_3_io_q_vk; 
  wire  FFs_3_io_q_busy; 
  wire [19:0] FFs_3_io_d_op; 
  wire [4:0] FFs_3_io_d_dest; 
  wire [4:0] FFs_3_io_d_qj; 
  wire [4:0] FFs_3_io_d_qk; 
  wire [31:0] FFs_3_io_d_a; 
  wire [31:0] FFs_3_io_d_vj; 
  wire [31:0] FFs_3_io_d_vk; 
  wire  FFs_3_io_d_busy; 
  wire  FFs_3_io_clear; 
  wire [1:0] _io_full_T_1 = h_ptr_io_q + 2'h1; 
  wire [31:0] FFs_io_0_q_vk = FFs_0_io_q_vk; 
  wire  FFs_io_0_q_busy = FFs_0_io_q_busy; 
  wire [31:0] FFs_io_0_q_a = FFs_0_io_q_a; 
  wire [31:0] FFs_io_0_q_vj = FFs_0_io_q_vj; 
  wire [4:0] FFs_io_0_q_qj = FFs_0_io_q_qj; 
  wire [4:0] FFs_io_0_q_qk = FFs_0_io_q_qk; 
  wire [19:0] FFs_io_0_q_op = FFs_0_io_q_op; 
  wire [4:0] FFs_io_0_q_dest = FFs_0_io_q_dest; 
  wire [131:0] io_queue_data_lo_lo = {FFs_io_0_q_op,FFs_io_0_q_dest,FFs_io_0_q_qj,FFs_io_0_q_qk,FFs_io_0_q_a,
    FFs_io_0_q_vj,FFs_io_0_q_vk,FFs_io_0_q_busy}; 
  wire [31:0] FFs_io_1_q_vk = FFs_1_io_q_vk; 
  wire  FFs_io_1_q_busy = FFs_1_io_q_busy; 
  wire [31:0] FFs_io_1_q_a = FFs_1_io_q_a; 
  wire [31:0] FFs_io_1_q_vj = FFs_1_io_q_vj; 
  wire [4:0] FFs_io_1_q_qj = FFs_1_io_q_qj; 
  wire [4:0] FFs_io_1_q_qk = FFs_1_io_q_qk; 
  wire [19:0] FFs_io_1_q_op = FFs_1_io_q_op; 
  wire [4:0] FFs_io_1_q_dest = FFs_1_io_q_dest; 
  wire [263:0] io_queue_data_lo = {FFs_io_1_q_op,FFs_io_1_q_dest,FFs_io_1_q_qj,FFs_io_1_q_qk,FFs_io_1_q_a,FFs_io_1_q_vj,
    FFs_io_1_q_vk,FFs_io_1_q_busy,io_queue_data_lo_lo}; 
  wire [31:0] FFs_io_2_q_vk = FFs_2_io_q_vk; 
  wire  FFs_io_2_q_busy = FFs_2_io_q_busy; 
  wire [31:0] FFs_io_2_q_a = FFs_2_io_q_a; 
  wire [31:0] FFs_io_2_q_vj = FFs_2_io_q_vj; 
  wire [4:0] FFs_io_2_q_qj = FFs_2_io_q_qj; 
  wire [4:0] FFs_io_2_q_qk = FFs_2_io_q_qk; 
  wire [19:0] FFs_io_2_q_op = FFs_2_io_q_op; 
  wire [4:0] FFs_io_2_q_dest = FFs_2_io_q_dest; 
  wire [131:0] io_queue_data_hi_lo = {FFs_io_2_q_op,FFs_io_2_q_dest,FFs_io_2_q_qj,FFs_io_2_q_qk,FFs_io_2_q_a,
    FFs_io_2_q_vj,FFs_io_2_q_vk,FFs_io_2_q_busy}; 
  wire [31:0] FFs_io_3_q_vk = FFs_3_io_q_vk; 
  wire  FFs_io_3_q_busy = FFs_3_io_q_busy; 
  wire [31:0] FFs_io_3_q_a = FFs_3_io_q_a; 
  wire [31:0] FFs_io_3_q_vj = FFs_3_io_q_vj; 
  wire [4:0] FFs_io_3_q_qj = FFs_3_io_q_qj; 
  wire [4:0] FFs_io_3_q_qk = FFs_3_io_q_qk; 
  wire [19:0] FFs_io_3_q_op = FFs_3_io_q_op; 
  wire [4:0] FFs_io_3_q_dest = FFs_3_io_q_dest; 
  wire [263:0] io_queue_data_hi = {FFs_io_3_q_op,FFs_io_3_q_dest,FFs_io_3_q_qj,FFs_io_3_q_qk,FFs_io_3_q_a,FFs_io_3_q_vj,
    FFs_io_3_q_vk,FFs_io_3_q_busy,io_queue_data_hi_lo}; 
  wire [31:0] _GEN_1 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_vk : FFs_io_0_q_vk; 
  wire [31:0] _GEN_2 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_vk : _GEN_1; 
  wire [31:0] _GEN_3 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_vk : _GEN_2; 
  wire  _GEN_5 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_busy : FFs_io_0_q_busy; 
  wire  _GEN_6 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_busy : _GEN_5; 
  wire  _GEN_7 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_busy : _GEN_6; 
  wire [31:0] _GEN_9 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_a : FFs_io_0_q_a; 
  wire [31:0] _GEN_10 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_a : _GEN_9; 
  wire [31:0] _GEN_11 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_a : _GEN_10; 
  wire [31:0] _GEN_13 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_vj : FFs_io_0_q_vj; 
  wire [31:0] _GEN_14 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_vj : _GEN_13; 
  wire [31:0] _GEN_15 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_vj : _GEN_14; 
  wire [96:0] io_deq_data_lo = {_GEN_11,_GEN_15,_GEN_3,_GEN_7}; 
  wire [4:0] _GEN_17 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_qj : FFs_io_0_q_qj; 
  wire [4:0] _GEN_18 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_qj : _GEN_17; 
  wire [4:0] _GEN_19 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_qj : _GEN_18; 
  wire [4:0] _GEN_21 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_qk : FFs_io_0_q_qk; 
  wire [4:0] _GEN_22 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_qk : _GEN_21; 
  wire [4:0] _GEN_23 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_qk : _GEN_22; 
  wire [19:0] _GEN_25 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_op : FFs_io_0_q_op; 
  wire [19:0] _GEN_26 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_op : _GEN_25; 
  wire [19:0] _GEN_27 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_op : _GEN_26; 
  wire [4:0] _GEN_29 = 2'h1 == t_ptr_io_q ? FFs_io_1_q_dest : FFs_io_0_q_dest; 
  wire [4:0] _GEN_30 = 2'h2 == t_ptr_io_q ? FFs_io_2_q_dest : _GEN_29; 
  wire [4:0] _GEN_31 = 2'h3 == t_ptr_io_q ? FFs_io_3_q_dest : _GEN_30; 
  wire [34:0] io_deq_data_hi = {_GEN_27,_GEN_31,_GEN_19,_GEN_23}; 
  wire  _T_1 = io_enq & ~io_full; 
  wire  _T_4 = io_deq & ~io_empty; 
  wire [1:0] _t_ptr_io_d_T_1 = t_ptr_io_q + 2'h1; 
  wire  _GEN_34 = io_update_entry[0] ? io_update_entry_data[0] : FFs_io_0_q_busy; 
  wire [31:0] _GEN_35 = io_update_entry[0] ? io_update_entry_data[32:1] : FFs_io_0_q_vk; 
  wire [31:0] _GEN_36 = io_update_entry[0] ? io_update_entry_data[64:33] : FFs_io_0_q_vj; 
  wire [31:0] _GEN_37 = io_update_entry[0] ? io_update_entry_data[96:65] : FFs_io_0_q_a; 
  wire [4:0] _GEN_38 = io_update_entry[0] ? io_update_entry_data[101:97] : FFs_io_0_q_qk; 
  wire [4:0] _GEN_39 = io_update_entry[0] ? io_update_entry_data[106:102] : FFs_io_0_q_qj; 
  wire [4:0] _GEN_40 = io_update_entry[0] ? io_update_entry_data[111:107] : FFs_io_0_q_dest; 
  wire [19:0] _GEN_41 = io_update_entry[0] ? io_update_entry_data[131:112] : FFs_io_0_q_op; 
  wire  _GEN_51 = io_update_entry[1] ? io_update_entry_data[132] : FFs_io_1_q_busy; 
  wire [31:0] _GEN_52 = io_update_entry[1] ? io_update_entry_data[164:133] : FFs_io_1_q_vk; 
  wire [31:0] _GEN_53 = io_update_entry[1] ? io_update_entry_data[196:165] : FFs_io_1_q_vj; 
  wire [31:0] _GEN_54 = io_update_entry[1] ? io_update_entry_data[228:197] : FFs_io_1_q_a; 
  wire [4:0] _GEN_55 = io_update_entry[1] ? io_update_entry_data[233:229] : FFs_io_1_q_qk; 
  wire [4:0] _GEN_56 = io_update_entry[1] ? io_update_entry_data[238:234] : FFs_io_1_q_qj; 
  wire [4:0] _GEN_57 = io_update_entry[1] ? io_update_entry_data[243:239] : FFs_io_1_q_dest; 
  wire [19:0] _GEN_58 = io_update_entry[1] ? io_update_entry_data[263:244] : FFs_io_1_q_op; 
  wire  _GEN_68 = io_update_entry[2] ? io_update_entry_data[264] : FFs_io_2_q_busy; 
  wire [31:0] _GEN_69 = io_update_entry[2] ? io_update_entry_data[296:265] : FFs_io_2_q_vk; 
  wire [31:0] _GEN_70 = io_update_entry[2] ? io_update_entry_data[328:297] : FFs_io_2_q_vj; 
  wire [31:0] _GEN_71 = io_update_entry[2] ? io_update_entry_data[360:329] : FFs_io_2_q_a; 
  wire [4:0] _GEN_72 = io_update_entry[2] ? io_update_entry_data[365:361] : FFs_io_2_q_qk; 
  wire [4:0] _GEN_73 = io_update_entry[2] ? io_update_entry_data[370:366] : FFs_io_2_q_qj; 
  wire [4:0] _GEN_74 = io_update_entry[2] ? io_update_entry_data[375:371] : FFs_io_2_q_dest; 
  wire [19:0] _GEN_75 = io_update_entry[2] ? io_update_entry_data[395:376] : FFs_io_2_q_op; 
  wire  _GEN_85 = io_update_entry[3] ? io_update_entry_data[396] : FFs_io_3_q_busy; 
  wire [31:0] _GEN_86 = io_update_entry[3] ? io_update_entry_data[428:397] : FFs_io_3_q_vk; 
  wire [31:0] _GEN_87 = io_update_entry[3] ? io_update_entry_data[460:429] : FFs_io_3_q_vj; 
  wire [31:0] _GEN_88 = io_update_entry[3] ? io_update_entry_data[492:461] : FFs_io_3_q_a; 
  wire [4:0] _GEN_89 = io_update_entry[3] ? io_update_entry_data[497:493] : FFs_io_3_q_qk; 
  wire [4:0] _GEN_90 = io_update_entry[3] ? io_update_entry_data[502:498] : FFs_io_3_q_qj; 
  wire [4:0] _GEN_91 = io_update_entry[3] ? io_update_entry_data[507:503] : FFs_io_3_q_dest; 
  wire [19:0] _GEN_92 = io_update_entry[3] ? io_update_entry_data[527:508] : FFs_io_3_q_op; 
  prim_ff_cl_5 h_ptr ( 
    .clock(h_ptr_clock),
    .reset(h_ptr_reset),
    .io_q(h_ptr_io_q),
    .io_d(h_ptr_io_d),
    .io_clear(h_ptr_io_clear)
  );
  prim_ff_cl_5 t_ptr ( 
    .clock(t_ptr_clock),
    .reset(t_ptr_reset),
    .io_q(t_ptr_io_q),
    .io_d(t_ptr_io_d),
    .io_clear(t_ptr_io_clear)
  );
  prim_ff_cl FFs_0 ( 
    .clock(FFs_0_clock),
    .reset(FFs_0_reset),
    .io_q_op(FFs_0_io_q_op),
    .io_q_dest(FFs_0_io_q_dest),
    .io_q_qj(FFs_0_io_q_qj),
    .io_q_qk(FFs_0_io_q_qk),
    .io_q_a(FFs_0_io_q_a),
    .io_q_vj(FFs_0_io_q_vj),
    .io_q_vk(FFs_0_io_q_vk),
    .io_q_busy(FFs_0_io_q_busy),
    .io_d_op(FFs_0_io_d_op),
    .io_d_dest(FFs_0_io_d_dest),
    .io_d_qj(FFs_0_io_d_qj),
    .io_d_qk(FFs_0_io_d_qk),
    .io_d_a(FFs_0_io_d_a),
    .io_d_vj(FFs_0_io_d_vj),
    .io_d_vk(FFs_0_io_d_vk),
    .io_d_busy(FFs_0_io_d_busy),
    .io_clear(FFs_0_io_clear)
  );
  prim_ff_cl FFs_1 ( 
    .clock(FFs_1_clock),
    .reset(FFs_1_reset),
    .io_q_op(FFs_1_io_q_op),
    .io_q_dest(FFs_1_io_q_dest),
    .io_q_qj(FFs_1_io_q_qj),
    .io_q_qk(FFs_1_io_q_qk),
    .io_q_a(FFs_1_io_q_a),
    .io_q_vj(FFs_1_io_q_vj),
    .io_q_vk(FFs_1_io_q_vk),
    .io_q_busy(FFs_1_io_q_busy),
    .io_d_op(FFs_1_io_d_op),
    .io_d_dest(FFs_1_io_d_dest),
    .io_d_qj(FFs_1_io_d_qj),
    .io_d_qk(FFs_1_io_d_qk),
    .io_d_a(FFs_1_io_d_a),
    .io_d_vj(FFs_1_io_d_vj),
    .io_d_vk(FFs_1_io_d_vk),
    .io_d_busy(FFs_1_io_d_busy),
    .io_clear(FFs_1_io_clear)
  );
  prim_ff_cl FFs_2 ( 
    .clock(FFs_2_clock),
    .reset(FFs_2_reset),
    .io_q_op(FFs_2_io_q_op),
    .io_q_dest(FFs_2_io_q_dest),
    .io_q_qj(FFs_2_io_q_qj),
    .io_q_qk(FFs_2_io_q_qk),
    .io_q_a(FFs_2_io_q_a),
    .io_q_vj(FFs_2_io_q_vj),
    .io_q_vk(FFs_2_io_q_vk),
    .io_q_busy(FFs_2_io_q_busy),
    .io_d_op(FFs_2_io_d_op),
    .io_d_dest(FFs_2_io_d_dest),
    .io_d_qj(FFs_2_io_d_qj),
    .io_d_qk(FFs_2_io_d_qk),
    .io_d_a(FFs_2_io_d_a),
    .io_d_vj(FFs_2_io_d_vj),
    .io_d_vk(FFs_2_io_d_vk),
    .io_d_busy(FFs_2_io_d_busy),
    .io_clear(FFs_2_io_clear)
  );
  prim_ff_cl FFs_3 ( 
    .clock(FFs_3_clock),
    .reset(FFs_3_reset),
    .io_q_op(FFs_3_io_q_op),
    .io_q_dest(FFs_3_io_q_dest),
    .io_q_qj(FFs_3_io_q_qj),
    .io_q_qk(FFs_3_io_q_qk),
    .io_q_a(FFs_3_io_q_a),
    .io_q_vj(FFs_3_io_q_vj),
    .io_q_vk(FFs_3_io_q_vk),
    .io_q_busy(FFs_3_io_q_busy),
    .io_d_op(FFs_3_io_d_op),
    .io_d_dest(FFs_3_io_d_dest),
    .io_d_qj(FFs_3_io_d_qj),
    .io_d_qk(FFs_3_io_d_qk),
    .io_d_a(FFs_3_io_d_a),
    .io_d_vj(FFs_3_io_d_vj),
    .io_d_vk(FFs_3_io_d_vk),
    .io_d_busy(FFs_3_io_d_busy),
    .io_clear(FFs_3_io_clear)
  );
  assign io_enq_idx = h_ptr_io_q; 
  assign io_deq_data = {io_deq_data_hi,io_deq_data_lo}; 
  assign io_deq_idx = t_ptr_io_q; 
  assign io_empty = h_ptr_io_q == t_ptr_io_q; 
  assign io_full = _io_full_T_1 == t_ptr_io_q; 
  assign io_queue_data = {io_queue_data_hi,io_queue_data_lo}; 
  assign h_ptr_clock = clock;
  assign h_ptr_reset = reset;
  assign h_ptr_io_d = io_enq & ~io_full ? _io_full_T_1 : h_ptr_io_q; 
  assign h_ptr_io_clear = io_clear; 
  assign t_ptr_clock = clock;
  assign t_ptr_reset = reset;
  assign t_ptr_io_d = io_deq & ~io_empty ? _t_ptr_io_d_T_1 : t_ptr_io_q; 
  assign t_ptr_io_clear = io_clear; 
  assign FFs_0_clock = clock;
  assign FFs_0_reset = reset;
  assign FFs_0_io_d_op = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[131:112] : _GEN_41; 
  assign FFs_0_io_d_dest = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[111:107] : _GEN_40; 
  assign FFs_0_io_d_qj = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[106:102] : _GEN_39; 
  assign FFs_0_io_d_qk = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[101:97] : _GEN_38; 
  assign FFs_0_io_d_a = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[96:65] : _GEN_37; 
  assign FFs_0_io_d_vj = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_36; 
  assign FFs_0_io_d_vk = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_35; 
  assign FFs_0_io_d_busy = 2'h0 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_34; 
  assign FFs_0_io_clear = 2'h0 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_1_clock = clock;
  assign FFs_1_reset = reset;
  assign FFs_1_io_d_op = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[131:112] : _GEN_58; 
  assign FFs_1_io_d_dest = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[111:107] : _GEN_57; 
  assign FFs_1_io_d_qj = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[106:102] : _GEN_56; 
  assign FFs_1_io_d_qk = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[101:97] : _GEN_55; 
  assign FFs_1_io_d_a = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[96:65] : _GEN_54; 
  assign FFs_1_io_d_vj = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_53; 
  assign FFs_1_io_d_vk = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_52; 
  assign FFs_1_io_d_busy = 2'h1 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_51; 
  assign FFs_1_io_clear = 2'h1 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_2_clock = clock;
  assign FFs_2_reset = reset;
  assign FFs_2_io_d_op = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[131:112] : _GEN_75; 
  assign FFs_2_io_d_dest = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[111:107] : _GEN_74; 
  assign FFs_2_io_d_qj = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[106:102] : _GEN_73; 
  assign FFs_2_io_d_qk = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[101:97] : _GEN_72; 
  assign FFs_2_io_d_a = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[96:65] : _GEN_71; 
  assign FFs_2_io_d_vj = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_70; 
  assign FFs_2_io_d_vk = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_69; 
  assign FFs_2_io_d_busy = 2'h2 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_68; 
  assign FFs_2_io_clear = 2'h2 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_3_clock = clock;
  assign FFs_3_reset = reset;
  assign FFs_3_io_d_op = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[131:112] : _GEN_92; 
  assign FFs_3_io_d_dest = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[111:107] : _GEN_91; 
  assign FFs_3_io_d_qj = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[106:102] : _GEN_90; 
  assign FFs_3_io_d_qk = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[101:97] : _GEN_89; 
  assign FFs_3_io_d_a = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[96:65] : _GEN_88; 
  assign FFs_3_io_d_vj = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_87; 
  assign FFs_3_io_d_vk = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_86; 
  assign FFs_3_io_d_busy = 2'h3 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_85; 
  assign FFs_3_io_clear = 2'h3 == io_deq_idx & _T_4 | io_clear; 
endmodule
module prim_ff_cl_17(
  input        clock,
  input        reset,
  output [3:0] io_q, 
  input  [3:0] io_d, 
  input        io_clear 
);
  reg [3:0] m_reg; 
  assign io_q = m_reg; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg <= 4'h0; 
    end else if (io_clear) begin 
      m_reg <= 4'h0;
    end else begin
      m_reg <= io_d;
    end
  end
endmodule
module prim_ff_cl_19(
  input         clock,
  input         reset,
  output [1:0]  io_q_rob_type, 
  output [31:0] io_q_rob_dest, 
  output [31:0] io_q_rob_value, 
  output        io_q_rob_ready, 
  input  [1:0]  io_d_rob_type, 
  input  [31:0] io_d_rob_dest, 
  input  [31:0] io_d_rob_value, 
  input         io_d_rob_ready, 
  input         io_clear 
);
  reg [1:0] m_reg_rob_type; 
  reg [31:0] m_reg_rob_dest; 
  reg [31:0] m_reg_rob_value; 
  reg  m_reg_rob_ready; 
  assign io_q_rob_type = m_reg_rob_type; 
  assign io_q_rob_dest = m_reg_rob_dest; 
  assign io_q_rob_value = m_reg_rob_value; 
  assign io_q_rob_ready = m_reg_rob_ready; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_rob_type <= 2'h0; 
    end else if (io_clear) begin 
      m_reg_rob_type <= 2'h0;
    end else begin
      m_reg_rob_type <= io_d_rob_type;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_rob_dest <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_rob_dest <= 32'h0;
    end else begin
      m_reg_rob_dest <= io_d_rob_dest;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_rob_value <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_rob_value <= 32'h0;
    end else begin
      m_reg_rob_value <= io_d_rob_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_rob_ready <= 1'h0; 
    end else if (io_clear) begin 
      m_reg_rob_ready <= 1'h0;
    end else begin
      m_reg_rob_ready <= io_d_rob_ready;
    end
  end
endmodule
module FIFO_2(
  input           clock,
  input           reset,
  input           io_clear, 
  input           io_enq, 
  input  [66:0]   io_enq_data, 
  output [3:0]    io_enq_idx, 
  input           io_deq, 
  output [66:0]   io_deq_data, 
  output [3:0]    io_deq_idx, 
  output          io_empty, 
  output          io_full, 
  output [1071:0] io_queue_data, 
  input  [15:0]   io_update_entry, 
  input  [1071:0] io_update_entry_data 
);
  wire  h_ptr_clock; 
  wire  h_ptr_reset; 
  wire [3:0] h_ptr_io_q; 
  wire [3:0] h_ptr_io_d; 
  wire  h_ptr_io_clear; 
  wire  t_ptr_clock; 
  wire  t_ptr_reset; 
  wire [3:0] t_ptr_io_q; 
  wire [3:0] t_ptr_io_d; 
  wire  t_ptr_io_clear; 
  wire  FFs_0_clock; 
  wire  FFs_0_reset; 
  wire [1:0] FFs_0_io_q_rob_type; 
  wire [31:0] FFs_0_io_q_rob_dest; 
  wire [31:0] FFs_0_io_q_rob_value; 
  wire  FFs_0_io_q_rob_ready; 
  wire [1:0] FFs_0_io_d_rob_type; 
  wire [31:0] FFs_0_io_d_rob_dest; 
  wire [31:0] FFs_0_io_d_rob_value; 
  wire  FFs_0_io_d_rob_ready; 
  wire  FFs_0_io_clear; 
  wire  FFs_1_clock; 
  wire  FFs_1_reset; 
  wire [1:0] FFs_1_io_q_rob_type; 
  wire [31:0] FFs_1_io_q_rob_dest; 
  wire [31:0] FFs_1_io_q_rob_value; 
  wire  FFs_1_io_q_rob_ready; 
  wire [1:0] FFs_1_io_d_rob_type; 
  wire [31:0] FFs_1_io_d_rob_dest; 
  wire [31:0] FFs_1_io_d_rob_value; 
  wire  FFs_1_io_d_rob_ready; 
  wire  FFs_1_io_clear; 
  wire  FFs_2_clock; 
  wire  FFs_2_reset; 
  wire [1:0] FFs_2_io_q_rob_type; 
  wire [31:0] FFs_2_io_q_rob_dest; 
  wire [31:0] FFs_2_io_q_rob_value; 
  wire  FFs_2_io_q_rob_ready; 
  wire [1:0] FFs_2_io_d_rob_type; 
  wire [31:0] FFs_2_io_d_rob_dest; 
  wire [31:0] FFs_2_io_d_rob_value; 
  wire  FFs_2_io_d_rob_ready; 
  wire  FFs_2_io_clear; 
  wire  FFs_3_clock; 
  wire  FFs_3_reset; 
  wire [1:0] FFs_3_io_q_rob_type; 
  wire [31:0] FFs_3_io_q_rob_dest; 
  wire [31:0] FFs_3_io_q_rob_value; 
  wire  FFs_3_io_q_rob_ready; 
  wire [1:0] FFs_3_io_d_rob_type; 
  wire [31:0] FFs_3_io_d_rob_dest; 
  wire [31:0] FFs_3_io_d_rob_value; 
  wire  FFs_3_io_d_rob_ready; 
  wire  FFs_3_io_clear; 
  wire  FFs_4_clock; 
  wire  FFs_4_reset; 
  wire [1:0] FFs_4_io_q_rob_type; 
  wire [31:0] FFs_4_io_q_rob_dest; 
  wire [31:0] FFs_4_io_q_rob_value; 
  wire  FFs_4_io_q_rob_ready; 
  wire [1:0] FFs_4_io_d_rob_type; 
  wire [31:0] FFs_4_io_d_rob_dest; 
  wire [31:0] FFs_4_io_d_rob_value; 
  wire  FFs_4_io_d_rob_ready; 
  wire  FFs_4_io_clear; 
  wire  FFs_5_clock; 
  wire  FFs_5_reset; 
  wire [1:0] FFs_5_io_q_rob_type; 
  wire [31:0] FFs_5_io_q_rob_dest; 
  wire [31:0] FFs_5_io_q_rob_value; 
  wire  FFs_5_io_q_rob_ready; 
  wire [1:0] FFs_5_io_d_rob_type; 
  wire [31:0] FFs_5_io_d_rob_dest; 
  wire [31:0] FFs_5_io_d_rob_value; 
  wire  FFs_5_io_d_rob_ready; 
  wire  FFs_5_io_clear; 
  wire  FFs_6_clock; 
  wire  FFs_6_reset; 
  wire [1:0] FFs_6_io_q_rob_type; 
  wire [31:0] FFs_6_io_q_rob_dest; 
  wire [31:0] FFs_6_io_q_rob_value; 
  wire  FFs_6_io_q_rob_ready; 
  wire [1:0] FFs_6_io_d_rob_type; 
  wire [31:0] FFs_6_io_d_rob_dest; 
  wire [31:0] FFs_6_io_d_rob_value; 
  wire  FFs_6_io_d_rob_ready; 
  wire  FFs_6_io_clear; 
  wire  FFs_7_clock; 
  wire  FFs_7_reset; 
  wire [1:0] FFs_7_io_q_rob_type; 
  wire [31:0] FFs_7_io_q_rob_dest; 
  wire [31:0] FFs_7_io_q_rob_value; 
  wire  FFs_7_io_q_rob_ready; 
  wire [1:0] FFs_7_io_d_rob_type; 
  wire [31:0] FFs_7_io_d_rob_dest; 
  wire [31:0] FFs_7_io_d_rob_value; 
  wire  FFs_7_io_d_rob_ready; 
  wire  FFs_7_io_clear; 
  wire  FFs_8_clock; 
  wire  FFs_8_reset; 
  wire [1:0] FFs_8_io_q_rob_type; 
  wire [31:0] FFs_8_io_q_rob_dest; 
  wire [31:0] FFs_8_io_q_rob_value; 
  wire  FFs_8_io_q_rob_ready; 
  wire [1:0] FFs_8_io_d_rob_type; 
  wire [31:0] FFs_8_io_d_rob_dest; 
  wire [31:0] FFs_8_io_d_rob_value; 
  wire  FFs_8_io_d_rob_ready; 
  wire  FFs_8_io_clear; 
  wire  FFs_9_clock; 
  wire  FFs_9_reset; 
  wire [1:0] FFs_9_io_q_rob_type; 
  wire [31:0] FFs_9_io_q_rob_dest; 
  wire [31:0] FFs_9_io_q_rob_value; 
  wire  FFs_9_io_q_rob_ready; 
  wire [1:0] FFs_9_io_d_rob_type; 
  wire [31:0] FFs_9_io_d_rob_dest; 
  wire [31:0] FFs_9_io_d_rob_value; 
  wire  FFs_9_io_d_rob_ready; 
  wire  FFs_9_io_clear; 
  wire  FFs_10_clock; 
  wire  FFs_10_reset; 
  wire [1:0] FFs_10_io_q_rob_type; 
  wire [31:0] FFs_10_io_q_rob_dest; 
  wire [31:0] FFs_10_io_q_rob_value; 
  wire  FFs_10_io_q_rob_ready; 
  wire [1:0] FFs_10_io_d_rob_type; 
  wire [31:0] FFs_10_io_d_rob_dest; 
  wire [31:0] FFs_10_io_d_rob_value; 
  wire  FFs_10_io_d_rob_ready; 
  wire  FFs_10_io_clear; 
  wire  FFs_11_clock; 
  wire  FFs_11_reset; 
  wire [1:0] FFs_11_io_q_rob_type; 
  wire [31:0] FFs_11_io_q_rob_dest; 
  wire [31:0] FFs_11_io_q_rob_value; 
  wire  FFs_11_io_q_rob_ready; 
  wire [1:0] FFs_11_io_d_rob_type; 
  wire [31:0] FFs_11_io_d_rob_dest; 
  wire [31:0] FFs_11_io_d_rob_value; 
  wire  FFs_11_io_d_rob_ready; 
  wire  FFs_11_io_clear; 
  wire  FFs_12_clock; 
  wire  FFs_12_reset; 
  wire [1:0] FFs_12_io_q_rob_type; 
  wire [31:0] FFs_12_io_q_rob_dest; 
  wire [31:0] FFs_12_io_q_rob_value; 
  wire  FFs_12_io_q_rob_ready; 
  wire [1:0] FFs_12_io_d_rob_type; 
  wire [31:0] FFs_12_io_d_rob_dest; 
  wire [31:0] FFs_12_io_d_rob_value; 
  wire  FFs_12_io_d_rob_ready; 
  wire  FFs_12_io_clear; 
  wire  FFs_13_clock; 
  wire  FFs_13_reset; 
  wire [1:0] FFs_13_io_q_rob_type; 
  wire [31:0] FFs_13_io_q_rob_dest; 
  wire [31:0] FFs_13_io_q_rob_value; 
  wire  FFs_13_io_q_rob_ready; 
  wire [1:0] FFs_13_io_d_rob_type; 
  wire [31:0] FFs_13_io_d_rob_dest; 
  wire [31:0] FFs_13_io_d_rob_value; 
  wire  FFs_13_io_d_rob_ready; 
  wire  FFs_13_io_clear; 
  wire  FFs_14_clock; 
  wire  FFs_14_reset; 
  wire [1:0] FFs_14_io_q_rob_type; 
  wire [31:0] FFs_14_io_q_rob_dest; 
  wire [31:0] FFs_14_io_q_rob_value; 
  wire  FFs_14_io_q_rob_ready; 
  wire [1:0] FFs_14_io_d_rob_type; 
  wire [31:0] FFs_14_io_d_rob_dest; 
  wire [31:0] FFs_14_io_d_rob_value; 
  wire  FFs_14_io_d_rob_ready; 
  wire  FFs_14_io_clear; 
  wire  FFs_15_clock; 
  wire  FFs_15_reset; 
  wire [1:0] FFs_15_io_q_rob_type; 
  wire [31:0] FFs_15_io_q_rob_dest; 
  wire [31:0] FFs_15_io_q_rob_value; 
  wire  FFs_15_io_q_rob_ready; 
  wire [1:0] FFs_15_io_d_rob_type; 
  wire [31:0] FFs_15_io_d_rob_dest; 
  wire [31:0] FFs_15_io_d_rob_value; 
  wire  FFs_15_io_d_rob_ready; 
  wire  FFs_15_io_clear; 
  wire [3:0] _io_full_T_1 = h_ptr_io_q + 4'h1; 
  wire [31:0] FFs_io_0_q_rob_value = FFs_0_io_q_rob_value; 
  wire  FFs_io_0_q_rob_ready = FFs_0_io_q_rob_ready; 
  wire [1:0] FFs_io_0_q_rob_type = FFs_0_io_q_rob_type; 
  wire [31:0] FFs_io_0_q_rob_dest = FFs_0_io_q_rob_dest; 
  wire [31:0] FFs_io_1_q_rob_value = FFs_1_io_q_rob_value; 
  wire  FFs_io_1_q_rob_ready = FFs_1_io_q_rob_ready; 
  wire [1:0] FFs_io_1_q_rob_type = FFs_1_io_q_rob_type; 
  wire [31:0] FFs_io_1_q_rob_dest = FFs_1_io_q_rob_dest; 
  wire [133:0] io_queue_data_lo_lo_lo = {FFs_io_1_q_rob_type,FFs_io_1_q_rob_dest,FFs_io_1_q_rob_value,
    FFs_io_1_q_rob_ready,FFs_io_0_q_rob_type,FFs_io_0_q_rob_dest,FFs_io_0_q_rob_value,FFs_io_0_q_rob_ready}; 
  wire [31:0] FFs_io_2_q_rob_value = FFs_2_io_q_rob_value; 
  wire  FFs_io_2_q_rob_ready = FFs_2_io_q_rob_ready; 
  wire [1:0] FFs_io_2_q_rob_type = FFs_2_io_q_rob_type; 
  wire [31:0] FFs_io_2_q_rob_dest = FFs_2_io_q_rob_dest; 
  wire [31:0] FFs_io_3_q_rob_value = FFs_3_io_q_rob_value; 
  wire  FFs_io_3_q_rob_ready = FFs_3_io_q_rob_ready; 
  wire [1:0] FFs_io_3_q_rob_type = FFs_3_io_q_rob_type; 
  wire [31:0] FFs_io_3_q_rob_dest = FFs_3_io_q_rob_dest; 
  wire [267:0] io_queue_data_lo_lo = {FFs_io_3_q_rob_type,FFs_io_3_q_rob_dest,FFs_io_3_q_rob_value,FFs_io_3_q_rob_ready,
    FFs_io_2_q_rob_type,FFs_io_2_q_rob_dest,FFs_io_2_q_rob_value,FFs_io_2_q_rob_ready,io_queue_data_lo_lo_lo}; 
  wire [31:0] FFs_io_4_q_rob_value = FFs_4_io_q_rob_value; 
  wire  FFs_io_4_q_rob_ready = FFs_4_io_q_rob_ready; 
  wire [1:0] FFs_io_4_q_rob_type = FFs_4_io_q_rob_type; 
  wire [31:0] FFs_io_4_q_rob_dest = FFs_4_io_q_rob_dest; 
  wire [31:0] FFs_io_5_q_rob_value = FFs_5_io_q_rob_value; 
  wire  FFs_io_5_q_rob_ready = FFs_5_io_q_rob_ready; 
  wire [1:0] FFs_io_5_q_rob_type = FFs_5_io_q_rob_type; 
  wire [31:0] FFs_io_5_q_rob_dest = FFs_5_io_q_rob_dest; 
  wire [133:0] io_queue_data_lo_hi_lo = {FFs_io_5_q_rob_type,FFs_io_5_q_rob_dest,FFs_io_5_q_rob_value,
    FFs_io_5_q_rob_ready,FFs_io_4_q_rob_type,FFs_io_4_q_rob_dest,FFs_io_4_q_rob_value,FFs_io_4_q_rob_ready}; 
  wire [31:0] FFs_io_6_q_rob_value = FFs_6_io_q_rob_value; 
  wire  FFs_io_6_q_rob_ready = FFs_6_io_q_rob_ready; 
  wire [1:0] FFs_io_6_q_rob_type = FFs_6_io_q_rob_type; 
  wire [31:0] FFs_io_6_q_rob_dest = FFs_6_io_q_rob_dest; 
  wire [31:0] FFs_io_7_q_rob_value = FFs_7_io_q_rob_value; 
  wire  FFs_io_7_q_rob_ready = FFs_7_io_q_rob_ready; 
  wire [1:0] FFs_io_7_q_rob_type = FFs_7_io_q_rob_type; 
  wire [31:0] FFs_io_7_q_rob_dest = FFs_7_io_q_rob_dest; 
  wire [535:0] io_queue_data_lo = {FFs_io_7_q_rob_type,FFs_io_7_q_rob_dest,FFs_io_7_q_rob_value,FFs_io_7_q_rob_ready,
    FFs_io_6_q_rob_type,FFs_io_6_q_rob_dest,FFs_io_6_q_rob_value,FFs_io_6_q_rob_ready,io_queue_data_lo_hi_lo,
    io_queue_data_lo_lo}; 
  wire [31:0] FFs_io_8_q_rob_value = FFs_8_io_q_rob_value; 
  wire  FFs_io_8_q_rob_ready = FFs_8_io_q_rob_ready; 
  wire [1:0] FFs_io_8_q_rob_type = FFs_8_io_q_rob_type; 
  wire [31:0] FFs_io_8_q_rob_dest = FFs_8_io_q_rob_dest; 
  wire [31:0] FFs_io_9_q_rob_value = FFs_9_io_q_rob_value; 
  wire  FFs_io_9_q_rob_ready = FFs_9_io_q_rob_ready; 
  wire [1:0] FFs_io_9_q_rob_type = FFs_9_io_q_rob_type; 
  wire [31:0] FFs_io_9_q_rob_dest = FFs_9_io_q_rob_dest; 
  wire [133:0] io_queue_data_hi_lo_lo = {FFs_io_9_q_rob_type,FFs_io_9_q_rob_dest,FFs_io_9_q_rob_value,
    FFs_io_9_q_rob_ready,FFs_io_8_q_rob_type,FFs_io_8_q_rob_dest,FFs_io_8_q_rob_value,FFs_io_8_q_rob_ready}; 
  wire [31:0] FFs_io_10_q_rob_value = FFs_10_io_q_rob_value; 
  wire  FFs_io_10_q_rob_ready = FFs_10_io_q_rob_ready; 
  wire [1:0] FFs_io_10_q_rob_type = FFs_10_io_q_rob_type; 
  wire [31:0] FFs_io_10_q_rob_dest = FFs_10_io_q_rob_dest; 
  wire [31:0] FFs_io_11_q_rob_value = FFs_11_io_q_rob_value; 
  wire  FFs_io_11_q_rob_ready = FFs_11_io_q_rob_ready; 
  wire [1:0] FFs_io_11_q_rob_type = FFs_11_io_q_rob_type; 
  wire [31:0] FFs_io_11_q_rob_dest = FFs_11_io_q_rob_dest; 
  wire [267:0] io_queue_data_hi_lo = {FFs_io_11_q_rob_type,FFs_io_11_q_rob_dest,FFs_io_11_q_rob_value,
    FFs_io_11_q_rob_ready,FFs_io_10_q_rob_type,FFs_io_10_q_rob_dest,FFs_io_10_q_rob_value,FFs_io_10_q_rob_ready,
    io_queue_data_hi_lo_lo}; 
  wire [31:0] FFs_io_12_q_rob_value = FFs_12_io_q_rob_value; 
  wire  FFs_io_12_q_rob_ready = FFs_12_io_q_rob_ready; 
  wire [1:0] FFs_io_12_q_rob_type = FFs_12_io_q_rob_type; 
  wire [31:0] FFs_io_12_q_rob_dest = FFs_12_io_q_rob_dest; 
  wire [31:0] FFs_io_13_q_rob_value = FFs_13_io_q_rob_value; 
  wire  FFs_io_13_q_rob_ready = FFs_13_io_q_rob_ready; 
  wire [1:0] FFs_io_13_q_rob_type = FFs_13_io_q_rob_type; 
  wire [31:0] FFs_io_13_q_rob_dest = FFs_13_io_q_rob_dest; 
  wire [133:0] io_queue_data_hi_hi_lo = {FFs_io_13_q_rob_type,FFs_io_13_q_rob_dest,FFs_io_13_q_rob_value,
    FFs_io_13_q_rob_ready,FFs_io_12_q_rob_type,FFs_io_12_q_rob_dest,FFs_io_12_q_rob_value,FFs_io_12_q_rob_ready}; 
  wire [31:0] FFs_io_14_q_rob_value = FFs_14_io_q_rob_value; 
  wire  FFs_io_14_q_rob_ready = FFs_14_io_q_rob_ready; 
  wire [1:0] FFs_io_14_q_rob_type = FFs_14_io_q_rob_type; 
  wire [31:0] FFs_io_14_q_rob_dest = FFs_14_io_q_rob_dest; 
  wire [31:0] FFs_io_15_q_rob_value = FFs_15_io_q_rob_value; 
  wire  FFs_io_15_q_rob_ready = FFs_15_io_q_rob_ready; 
  wire [1:0] FFs_io_15_q_rob_type = FFs_15_io_q_rob_type; 
  wire [31:0] FFs_io_15_q_rob_dest = FFs_15_io_q_rob_dest; 
  wire [535:0] io_queue_data_hi = {FFs_io_15_q_rob_type,FFs_io_15_q_rob_dest,FFs_io_15_q_rob_value,FFs_io_15_q_rob_ready
    ,FFs_io_14_q_rob_type,FFs_io_14_q_rob_dest,FFs_io_14_q_rob_value,FFs_io_14_q_rob_ready,io_queue_data_hi_hi_lo,
    io_queue_data_hi_lo}; 
  wire [31:0] _GEN_1 = 4'h1 == t_ptr_io_q ? FFs_io_1_q_rob_value : FFs_io_0_q_rob_value; 
  wire [31:0] _GEN_2 = 4'h2 == t_ptr_io_q ? FFs_io_2_q_rob_value : _GEN_1; 
  wire [31:0] _GEN_3 = 4'h3 == t_ptr_io_q ? FFs_io_3_q_rob_value : _GEN_2; 
  wire [31:0] _GEN_4 = 4'h4 == t_ptr_io_q ? FFs_io_4_q_rob_value : _GEN_3; 
  wire [31:0] _GEN_5 = 4'h5 == t_ptr_io_q ? FFs_io_5_q_rob_value : _GEN_4; 
  wire [31:0] _GEN_6 = 4'h6 == t_ptr_io_q ? FFs_io_6_q_rob_value : _GEN_5; 
  wire [31:0] _GEN_7 = 4'h7 == t_ptr_io_q ? FFs_io_7_q_rob_value : _GEN_6; 
  wire [31:0] _GEN_8 = 4'h8 == t_ptr_io_q ? FFs_io_8_q_rob_value : _GEN_7; 
  wire [31:0] _GEN_9 = 4'h9 == t_ptr_io_q ? FFs_io_9_q_rob_value : _GEN_8; 
  wire [31:0] _GEN_10 = 4'ha == t_ptr_io_q ? FFs_io_10_q_rob_value : _GEN_9; 
  wire [31:0] _GEN_11 = 4'hb == t_ptr_io_q ? FFs_io_11_q_rob_value : _GEN_10; 
  wire [31:0] _GEN_12 = 4'hc == t_ptr_io_q ? FFs_io_12_q_rob_value : _GEN_11; 
  wire [31:0] _GEN_13 = 4'hd == t_ptr_io_q ? FFs_io_13_q_rob_value : _GEN_12; 
  wire [31:0] _GEN_14 = 4'he == t_ptr_io_q ? FFs_io_14_q_rob_value : _GEN_13; 
  wire [31:0] _GEN_15 = 4'hf == t_ptr_io_q ? FFs_io_15_q_rob_value : _GEN_14; 
  wire  _GEN_17 = 4'h1 == t_ptr_io_q ? FFs_io_1_q_rob_ready : FFs_io_0_q_rob_ready; 
  wire  _GEN_18 = 4'h2 == t_ptr_io_q ? FFs_io_2_q_rob_ready : _GEN_17; 
  wire  _GEN_19 = 4'h3 == t_ptr_io_q ? FFs_io_3_q_rob_ready : _GEN_18; 
  wire  _GEN_20 = 4'h4 == t_ptr_io_q ? FFs_io_4_q_rob_ready : _GEN_19; 
  wire  _GEN_21 = 4'h5 == t_ptr_io_q ? FFs_io_5_q_rob_ready : _GEN_20; 
  wire  _GEN_22 = 4'h6 == t_ptr_io_q ? FFs_io_6_q_rob_ready : _GEN_21; 
  wire  _GEN_23 = 4'h7 == t_ptr_io_q ? FFs_io_7_q_rob_ready : _GEN_22; 
  wire  _GEN_24 = 4'h8 == t_ptr_io_q ? FFs_io_8_q_rob_ready : _GEN_23; 
  wire  _GEN_25 = 4'h9 == t_ptr_io_q ? FFs_io_9_q_rob_ready : _GEN_24; 
  wire  _GEN_26 = 4'ha == t_ptr_io_q ? FFs_io_10_q_rob_ready : _GEN_25; 
  wire  _GEN_27 = 4'hb == t_ptr_io_q ? FFs_io_11_q_rob_ready : _GEN_26; 
  wire  _GEN_28 = 4'hc == t_ptr_io_q ? FFs_io_12_q_rob_ready : _GEN_27; 
  wire  _GEN_29 = 4'hd == t_ptr_io_q ? FFs_io_13_q_rob_ready : _GEN_28; 
  wire  _GEN_30 = 4'he == t_ptr_io_q ? FFs_io_14_q_rob_ready : _GEN_29; 
  wire  _GEN_31 = 4'hf == t_ptr_io_q ? FFs_io_15_q_rob_ready : _GEN_30; 
  wire [32:0] io_deq_data_lo = {_GEN_15,_GEN_31}; 
  wire [1:0] _GEN_33 = 4'h1 == t_ptr_io_q ? FFs_io_1_q_rob_type : FFs_io_0_q_rob_type; 
  wire [1:0] _GEN_34 = 4'h2 == t_ptr_io_q ? FFs_io_2_q_rob_type : _GEN_33; 
  wire [1:0] _GEN_35 = 4'h3 == t_ptr_io_q ? FFs_io_3_q_rob_type : _GEN_34; 
  wire [1:0] _GEN_36 = 4'h4 == t_ptr_io_q ? FFs_io_4_q_rob_type : _GEN_35; 
  wire [1:0] _GEN_37 = 4'h5 == t_ptr_io_q ? FFs_io_5_q_rob_type : _GEN_36; 
  wire [1:0] _GEN_38 = 4'h6 == t_ptr_io_q ? FFs_io_6_q_rob_type : _GEN_37; 
  wire [1:0] _GEN_39 = 4'h7 == t_ptr_io_q ? FFs_io_7_q_rob_type : _GEN_38; 
  wire [1:0] _GEN_40 = 4'h8 == t_ptr_io_q ? FFs_io_8_q_rob_type : _GEN_39; 
  wire [1:0] _GEN_41 = 4'h9 == t_ptr_io_q ? FFs_io_9_q_rob_type : _GEN_40; 
  wire [1:0] _GEN_42 = 4'ha == t_ptr_io_q ? FFs_io_10_q_rob_type : _GEN_41; 
  wire [1:0] _GEN_43 = 4'hb == t_ptr_io_q ? FFs_io_11_q_rob_type : _GEN_42; 
  wire [1:0] _GEN_44 = 4'hc == t_ptr_io_q ? FFs_io_12_q_rob_type : _GEN_43; 
  wire [1:0] _GEN_45 = 4'hd == t_ptr_io_q ? FFs_io_13_q_rob_type : _GEN_44; 
  wire [1:0] _GEN_46 = 4'he == t_ptr_io_q ? FFs_io_14_q_rob_type : _GEN_45; 
  wire [1:0] _GEN_47 = 4'hf == t_ptr_io_q ? FFs_io_15_q_rob_type : _GEN_46; 
  wire [31:0] _GEN_49 = 4'h1 == t_ptr_io_q ? FFs_io_1_q_rob_dest : FFs_io_0_q_rob_dest; 
  wire [31:0] _GEN_50 = 4'h2 == t_ptr_io_q ? FFs_io_2_q_rob_dest : _GEN_49; 
  wire [31:0] _GEN_51 = 4'h3 == t_ptr_io_q ? FFs_io_3_q_rob_dest : _GEN_50; 
  wire [31:0] _GEN_52 = 4'h4 == t_ptr_io_q ? FFs_io_4_q_rob_dest : _GEN_51; 
  wire [31:0] _GEN_53 = 4'h5 == t_ptr_io_q ? FFs_io_5_q_rob_dest : _GEN_52; 
  wire [31:0] _GEN_54 = 4'h6 == t_ptr_io_q ? FFs_io_6_q_rob_dest : _GEN_53; 
  wire [31:0] _GEN_55 = 4'h7 == t_ptr_io_q ? FFs_io_7_q_rob_dest : _GEN_54; 
  wire [31:0] _GEN_56 = 4'h8 == t_ptr_io_q ? FFs_io_8_q_rob_dest : _GEN_55; 
  wire [31:0] _GEN_57 = 4'h9 == t_ptr_io_q ? FFs_io_9_q_rob_dest : _GEN_56; 
  wire [31:0] _GEN_58 = 4'ha == t_ptr_io_q ? FFs_io_10_q_rob_dest : _GEN_57; 
  wire [31:0] _GEN_59 = 4'hb == t_ptr_io_q ? FFs_io_11_q_rob_dest : _GEN_58; 
  wire [31:0] _GEN_60 = 4'hc == t_ptr_io_q ? FFs_io_12_q_rob_dest : _GEN_59; 
  wire [31:0] _GEN_61 = 4'hd == t_ptr_io_q ? FFs_io_13_q_rob_dest : _GEN_60; 
  wire [31:0] _GEN_62 = 4'he == t_ptr_io_q ? FFs_io_14_q_rob_dest : _GEN_61; 
  wire [31:0] _GEN_63 = 4'hf == t_ptr_io_q ? FFs_io_15_q_rob_dest : _GEN_62; 
  wire [33:0] io_deq_data_hi = {_GEN_47,_GEN_63}; 
  wire  _T_1 = io_enq & ~io_full; 
  wire  _T_4 = io_deq & ~io_empty; 
  wire [3:0] _t_ptr_io_d_T_1 = t_ptr_io_q + 4'h1; 
  wire  _GEN_66 = io_update_entry[0] ? io_update_entry_data[0] : FFs_io_0_q_rob_ready; 
  wire [31:0] _GEN_67 = io_update_entry[0] ? io_update_entry_data[32:1] : FFs_io_0_q_rob_value; 
  wire [31:0] _GEN_68 = io_update_entry[0] ? io_update_entry_data[64:33] : FFs_io_0_q_rob_dest; 
  wire [1:0] _GEN_69 = io_update_entry[0] ? io_update_entry_data[66:65] : FFs_io_0_q_rob_type; 
  wire  _GEN_75 = io_update_entry[1] ? io_update_entry_data[67] : FFs_io_1_q_rob_ready; 
  wire [31:0] _GEN_76 = io_update_entry[1] ? io_update_entry_data[99:68] : FFs_io_1_q_rob_value; 
  wire [31:0] _GEN_77 = io_update_entry[1] ? io_update_entry_data[131:100] : FFs_io_1_q_rob_dest; 
  wire [1:0] _GEN_78 = io_update_entry[1] ? io_update_entry_data[133:132] : FFs_io_1_q_rob_type; 
  wire  _GEN_84 = io_update_entry[2] ? io_update_entry_data[134] : FFs_io_2_q_rob_ready; 
  wire [31:0] _GEN_85 = io_update_entry[2] ? io_update_entry_data[166:135] : FFs_io_2_q_rob_value; 
  wire [31:0] _GEN_86 = io_update_entry[2] ? io_update_entry_data[198:167] : FFs_io_2_q_rob_dest; 
  wire [1:0] _GEN_87 = io_update_entry[2] ? io_update_entry_data[200:199] : FFs_io_2_q_rob_type; 
  wire  _GEN_93 = io_update_entry[3] ? io_update_entry_data[201] : FFs_io_3_q_rob_ready; 
  wire [31:0] _GEN_94 = io_update_entry[3] ? io_update_entry_data[233:202] : FFs_io_3_q_rob_value; 
  wire [31:0] _GEN_95 = io_update_entry[3] ? io_update_entry_data[265:234] : FFs_io_3_q_rob_dest; 
  wire [1:0] _GEN_96 = io_update_entry[3] ? io_update_entry_data[267:266] : FFs_io_3_q_rob_type; 
  wire  _GEN_102 = io_update_entry[4] ? io_update_entry_data[268] : FFs_io_4_q_rob_ready; 
  wire [31:0] _GEN_103 = io_update_entry[4] ? io_update_entry_data[300:269] : FFs_io_4_q_rob_value; 
  wire [31:0] _GEN_104 = io_update_entry[4] ? io_update_entry_data[332:301] : FFs_io_4_q_rob_dest; 
  wire [1:0] _GEN_105 = io_update_entry[4] ? io_update_entry_data[334:333] : FFs_io_4_q_rob_type; 
  wire  _GEN_111 = io_update_entry[5] ? io_update_entry_data[335] : FFs_io_5_q_rob_ready; 
  wire [31:0] _GEN_112 = io_update_entry[5] ? io_update_entry_data[367:336] : FFs_io_5_q_rob_value; 
  wire [31:0] _GEN_113 = io_update_entry[5] ? io_update_entry_data[399:368] : FFs_io_5_q_rob_dest; 
  wire [1:0] _GEN_114 = io_update_entry[5] ? io_update_entry_data[401:400] : FFs_io_5_q_rob_type; 
  wire  _GEN_120 = io_update_entry[6] ? io_update_entry_data[402] : FFs_io_6_q_rob_ready; 
  wire [31:0] _GEN_121 = io_update_entry[6] ? io_update_entry_data[434:403] : FFs_io_6_q_rob_value; 
  wire [31:0] _GEN_122 = io_update_entry[6] ? io_update_entry_data[466:435] : FFs_io_6_q_rob_dest; 
  wire [1:0] _GEN_123 = io_update_entry[6] ? io_update_entry_data[468:467] : FFs_io_6_q_rob_type; 
  wire  _GEN_129 = io_update_entry[7] ? io_update_entry_data[469] : FFs_io_7_q_rob_ready; 
  wire [31:0] _GEN_130 = io_update_entry[7] ? io_update_entry_data[501:470] : FFs_io_7_q_rob_value; 
  wire [31:0] _GEN_131 = io_update_entry[7] ? io_update_entry_data[533:502] : FFs_io_7_q_rob_dest; 
  wire [1:0] _GEN_132 = io_update_entry[7] ? io_update_entry_data[535:534] : FFs_io_7_q_rob_type; 
  wire  _GEN_138 = io_update_entry[8] ? io_update_entry_data[536] : FFs_io_8_q_rob_ready; 
  wire [31:0] _GEN_139 = io_update_entry[8] ? io_update_entry_data[568:537] : FFs_io_8_q_rob_value; 
  wire [31:0] _GEN_140 = io_update_entry[8] ? io_update_entry_data[600:569] : FFs_io_8_q_rob_dest; 
  wire [1:0] _GEN_141 = io_update_entry[8] ? io_update_entry_data[602:601] : FFs_io_8_q_rob_type; 
  wire  _GEN_147 = io_update_entry[9] ? io_update_entry_data[603] : FFs_io_9_q_rob_ready; 
  wire [31:0] _GEN_148 = io_update_entry[9] ? io_update_entry_data[635:604] : FFs_io_9_q_rob_value; 
  wire [31:0] _GEN_149 = io_update_entry[9] ? io_update_entry_data[667:636] : FFs_io_9_q_rob_dest; 
  wire [1:0] _GEN_150 = io_update_entry[9] ? io_update_entry_data[669:668] : FFs_io_9_q_rob_type; 
  wire  _GEN_156 = io_update_entry[10] ? io_update_entry_data[670] : FFs_io_10_q_rob_ready; 
  wire [31:0] _GEN_157 = io_update_entry[10] ? io_update_entry_data[702:671] : FFs_io_10_q_rob_value; 
  wire [31:0] _GEN_158 = io_update_entry[10] ? io_update_entry_data[734:703] : FFs_io_10_q_rob_dest; 
  wire [1:0] _GEN_159 = io_update_entry[10] ? io_update_entry_data[736:735] : FFs_io_10_q_rob_type; 
  wire  _GEN_165 = io_update_entry[11] ? io_update_entry_data[737] : FFs_io_11_q_rob_ready; 
  wire [31:0] _GEN_166 = io_update_entry[11] ? io_update_entry_data[769:738] : FFs_io_11_q_rob_value; 
  wire [31:0] _GEN_167 = io_update_entry[11] ? io_update_entry_data[801:770] : FFs_io_11_q_rob_dest; 
  wire [1:0] _GEN_168 = io_update_entry[11] ? io_update_entry_data[803:802] : FFs_io_11_q_rob_type; 
  wire  _GEN_174 = io_update_entry[12] ? io_update_entry_data[804] : FFs_io_12_q_rob_ready; 
  wire [31:0] _GEN_175 = io_update_entry[12] ? io_update_entry_data[836:805] : FFs_io_12_q_rob_value; 
  wire [31:0] _GEN_176 = io_update_entry[12] ? io_update_entry_data[868:837] : FFs_io_12_q_rob_dest; 
  wire [1:0] _GEN_177 = io_update_entry[12] ? io_update_entry_data[870:869] : FFs_io_12_q_rob_type; 
  wire  _GEN_183 = io_update_entry[13] ? io_update_entry_data[871] : FFs_io_13_q_rob_ready; 
  wire [31:0] _GEN_184 = io_update_entry[13] ? io_update_entry_data[903:872] : FFs_io_13_q_rob_value; 
  wire [31:0] _GEN_185 = io_update_entry[13] ? io_update_entry_data[935:904] : FFs_io_13_q_rob_dest; 
  wire [1:0] _GEN_186 = io_update_entry[13] ? io_update_entry_data[937:936] : FFs_io_13_q_rob_type; 
  wire  _GEN_192 = io_update_entry[14] ? io_update_entry_data[938] : FFs_io_14_q_rob_ready; 
  wire [31:0] _GEN_193 = io_update_entry[14] ? io_update_entry_data[970:939] : FFs_io_14_q_rob_value; 
  wire [31:0] _GEN_194 = io_update_entry[14] ? io_update_entry_data[1002:971] : FFs_io_14_q_rob_dest; 
  wire [1:0] _GEN_195 = io_update_entry[14] ? io_update_entry_data[1004:1003] : FFs_io_14_q_rob_type; 
  wire  _GEN_201 = io_update_entry[15] ? io_update_entry_data[1005] : FFs_io_15_q_rob_ready; 
  wire [31:0] _GEN_202 = io_update_entry[15] ? io_update_entry_data[1037:1006] : FFs_io_15_q_rob_value; 
  wire [31:0] _GEN_203 = io_update_entry[15] ? io_update_entry_data[1069:1038] : FFs_io_15_q_rob_dest; 
  wire [1:0] _GEN_204 = io_update_entry[15] ? io_update_entry_data[1071:1070] : FFs_io_15_q_rob_type; 
  prim_ff_cl_17 h_ptr ( 
    .clock(h_ptr_clock),
    .reset(h_ptr_reset),
    .io_q(h_ptr_io_q),
    .io_d(h_ptr_io_d),
    .io_clear(h_ptr_io_clear)
  );
  prim_ff_cl_17 t_ptr ( 
    .clock(t_ptr_clock),
    .reset(t_ptr_reset),
    .io_q(t_ptr_io_q),
    .io_d(t_ptr_io_d),
    .io_clear(t_ptr_io_clear)
  );
  prim_ff_cl_19 FFs_0 ( 
    .clock(FFs_0_clock),
    .reset(FFs_0_reset),
    .io_q_rob_type(FFs_0_io_q_rob_type),
    .io_q_rob_dest(FFs_0_io_q_rob_dest),
    .io_q_rob_value(FFs_0_io_q_rob_value),
    .io_q_rob_ready(FFs_0_io_q_rob_ready),
    .io_d_rob_type(FFs_0_io_d_rob_type),
    .io_d_rob_dest(FFs_0_io_d_rob_dest),
    .io_d_rob_value(FFs_0_io_d_rob_value),
    .io_d_rob_ready(FFs_0_io_d_rob_ready),
    .io_clear(FFs_0_io_clear)
  );
  prim_ff_cl_19 FFs_1 ( 
    .clock(FFs_1_clock),
    .reset(FFs_1_reset),
    .io_q_rob_type(FFs_1_io_q_rob_type),
    .io_q_rob_dest(FFs_1_io_q_rob_dest),
    .io_q_rob_value(FFs_1_io_q_rob_value),
    .io_q_rob_ready(FFs_1_io_q_rob_ready),
    .io_d_rob_type(FFs_1_io_d_rob_type),
    .io_d_rob_dest(FFs_1_io_d_rob_dest),
    .io_d_rob_value(FFs_1_io_d_rob_value),
    .io_d_rob_ready(FFs_1_io_d_rob_ready),
    .io_clear(FFs_1_io_clear)
  );
  prim_ff_cl_19 FFs_2 ( 
    .clock(FFs_2_clock),
    .reset(FFs_2_reset),
    .io_q_rob_type(FFs_2_io_q_rob_type),
    .io_q_rob_dest(FFs_2_io_q_rob_dest),
    .io_q_rob_value(FFs_2_io_q_rob_value),
    .io_q_rob_ready(FFs_2_io_q_rob_ready),
    .io_d_rob_type(FFs_2_io_d_rob_type),
    .io_d_rob_dest(FFs_2_io_d_rob_dest),
    .io_d_rob_value(FFs_2_io_d_rob_value),
    .io_d_rob_ready(FFs_2_io_d_rob_ready),
    .io_clear(FFs_2_io_clear)
  );
  prim_ff_cl_19 FFs_3 ( 
    .clock(FFs_3_clock),
    .reset(FFs_3_reset),
    .io_q_rob_type(FFs_3_io_q_rob_type),
    .io_q_rob_dest(FFs_3_io_q_rob_dest),
    .io_q_rob_value(FFs_3_io_q_rob_value),
    .io_q_rob_ready(FFs_3_io_q_rob_ready),
    .io_d_rob_type(FFs_3_io_d_rob_type),
    .io_d_rob_dest(FFs_3_io_d_rob_dest),
    .io_d_rob_value(FFs_3_io_d_rob_value),
    .io_d_rob_ready(FFs_3_io_d_rob_ready),
    .io_clear(FFs_3_io_clear)
  );
  prim_ff_cl_19 FFs_4 ( 
    .clock(FFs_4_clock),
    .reset(FFs_4_reset),
    .io_q_rob_type(FFs_4_io_q_rob_type),
    .io_q_rob_dest(FFs_4_io_q_rob_dest),
    .io_q_rob_value(FFs_4_io_q_rob_value),
    .io_q_rob_ready(FFs_4_io_q_rob_ready),
    .io_d_rob_type(FFs_4_io_d_rob_type),
    .io_d_rob_dest(FFs_4_io_d_rob_dest),
    .io_d_rob_value(FFs_4_io_d_rob_value),
    .io_d_rob_ready(FFs_4_io_d_rob_ready),
    .io_clear(FFs_4_io_clear)
  );
  prim_ff_cl_19 FFs_5 ( 
    .clock(FFs_5_clock),
    .reset(FFs_5_reset),
    .io_q_rob_type(FFs_5_io_q_rob_type),
    .io_q_rob_dest(FFs_5_io_q_rob_dest),
    .io_q_rob_value(FFs_5_io_q_rob_value),
    .io_q_rob_ready(FFs_5_io_q_rob_ready),
    .io_d_rob_type(FFs_5_io_d_rob_type),
    .io_d_rob_dest(FFs_5_io_d_rob_dest),
    .io_d_rob_value(FFs_5_io_d_rob_value),
    .io_d_rob_ready(FFs_5_io_d_rob_ready),
    .io_clear(FFs_5_io_clear)
  );
  prim_ff_cl_19 FFs_6 ( 
    .clock(FFs_6_clock),
    .reset(FFs_6_reset),
    .io_q_rob_type(FFs_6_io_q_rob_type),
    .io_q_rob_dest(FFs_6_io_q_rob_dest),
    .io_q_rob_value(FFs_6_io_q_rob_value),
    .io_q_rob_ready(FFs_6_io_q_rob_ready),
    .io_d_rob_type(FFs_6_io_d_rob_type),
    .io_d_rob_dest(FFs_6_io_d_rob_dest),
    .io_d_rob_value(FFs_6_io_d_rob_value),
    .io_d_rob_ready(FFs_6_io_d_rob_ready),
    .io_clear(FFs_6_io_clear)
  );
  prim_ff_cl_19 FFs_7 ( 
    .clock(FFs_7_clock),
    .reset(FFs_7_reset),
    .io_q_rob_type(FFs_7_io_q_rob_type),
    .io_q_rob_dest(FFs_7_io_q_rob_dest),
    .io_q_rob_value(FFs_7_io_q_rob_value),
    .io_q_rob_ready(FFs_7_io_q_rob_ready),
    .io_d_rob_type(FFs_7_io_d_rob_type),
    .io_d_rob_dest(FFs_7_io_d_rob_dest),
    .io_d_rob_value(FFs_7_io_d_rob_value),
    .io_d_rob_ready(FFs_7_io_d_rob_ready),
    .io_clear(FFs_7_io_clear)
  );
  prim_ff_cl_19 FFs_8 ( 
    .clock(FFs_8_clock),
    .reset(FFs_8_reset),
    .io_q_rob_type(FFs_8_io_q_rob_type),
    .io_q_rob_dest(FFs_8_io_q_rob_dest),
    .io_q_rob_value(FFs_8_io_q_rob_value),
    .io_q_rob_ready(FFs_8_io_q_rob_ready),
    .io_d_rob_type(FFs_8_io_d_rob_type),
    .io_d_rob_dest(FFs_8_io_d_rob_dest),
    .io_d_rob_value(FFs_8_io_d_rob_value),
    .io_d_rob_ready(FFs_8_io_d_rob_ready),
    .io_clear(FFs_8_io_clear)
  );
  prim_ff_cl_19 FFs_9 ( 
    .clock(FFs_9_clock),
    .reset(FFs_9_reset),
    .io_q_rob_type(FFs_9_io_q_rob_type),
    .io_q_rob_dest(FFs_9_io_q_rob_dest),
    .io_q_rob_value(FFs_9_io_q_rob_value),
    .io_q_rob_ready(FFs_9_io_q_rob_ready),
    .io_d_rob_type(FFs_9_io_d_rob_type),
    .io_d_rob_dest(FFs_9_io_d_rob_dest),
    .io_d_rob_value(FFs_9_io_d_rob_value),
    .io_d_rob_ready(FFs_9_io_d_rob_ready),
    .io_clear(FFs_9_io_clear)
  );
  prim_ff_cl_19 FFs_10 ( 
    .clock(FFs_10_clock),
    .reset(FFs_10_reset),
    .io_q_rob_type(FFs_10_io_q_rob_type),
    .io_q_rob_dest(FFs_10_io_q_rob_dest),
    .io_q_rob_value(FFs_10_io_q_rob_value),
    .io_q_rob_ready(FFs_10_io_q_rob_ready),
    .io_d_rob_type(FFs_10_io_d_rob_type),
    .io_d_rob_dest(FFs_10_io_d_rob_dest),
    .io_d_rob_value(FFs_10_io_d_rob_value),
    .io_d_rob_ready(FFs_10_io_d_rob_ready),
    .io_clear(FFs_10_io_clear)
  );
  prim_ff_cl_19 FFs_11 ( 
    .clock(FFs_11_clock),
    .reset(FFs_11_reset),
    .io_q_rob_type(FFs_11_io_q_rob_type),
    .io_q_rob_dest(FFs_11_io_q_rob_dest),
    .io_q_rob_value(FFs_11_io_q_rob_value),
    .io_q_rob_ready(FFs_11_io_q_rob_ready),
    .io_d_rob_type(FFs_11_io_d_rob_type),
    .io_d_rob_dest(FFs_11_io_d_rob_dest),
    .io_d_rob_value(FFs_11_io_d_rob_value),
    .io_d_rob_ready(FFs_11_io_d_rob_ready),
    .io_clear(FFs_11_io_clear)
  );
  prim_ff_cl_19 FFs_12 ( 
    .clock(FFs_12_clock),
    .reset(FFs_12_reset),
    .io_q_rob_type(FFs_12_io_q_rob_type),
    .io_q_rob_dest(FFs_12_io_q_rob_dest),
    .io_q_rob_value(FFs_12_io_q_rob_value),
    .io_q_rob_ready(FFs_12_io_q_rob_ready),
    .io_d_rob_type(FFs_12_io_d_rob_type),
    .io_d_rob_dest(FFs_12_io_d_rob_dest),
    .io_d_rob_value(FFs_12_io_d_rob_value),
    .io_d_rob_ready(FFs_12_io_d_rob_ready),
    .io_clear(FFs_12_io_clear)
  );
  prim_ff_cl_19 FFs_13 ( 
    .clock(FFs_13_clock),
    .reset(FFs_13_reset),
    .io_q_rob_type(FFs_13_io_q_rob_type),
    .io_q_rob_dest(FFs_13_io_q_rob_dest),
    .io_q_rob_value(FFs_13_io_q_rob_value),
    .io_q_rob_ready(FFs_13_io_q_rob_ready),
    .io_d_rob_type(FFs_13_io_d_rob_type),
    .io_d_rob_dest(FFs_13_io_d_rob_dest),
    .io_d_rob_value(FFs_13_io_d_rob_value),
    .io_d_rob_ready(FFs_13_io_d_rob_ready),
    .io_clear(FFs_13_io_clear)
  );
  prim_ff_cl_19 FFs_14 ( 
    .clock(FFs_14_clock),
    .reset(FFs_14_reset),
    .io_q_rob_type(FFs_14_io_q_rob_type),
    .io_q_rob_dest(FFs_14_io_q_rob_dest),
    .io_q_rob_value(FFs_14_io_q_rob_value),
    .io_q_rob_ready(FFs_14_io_q_rob_ready),
    .io_d_rob_type(FFs_14_io_d_rob_type),
    .io_d_rob_dest(FFs_14_io_d_rob_dest),
    .io_d_rob_value(FFs_14_io_d_rob_value),
    .io_d_rob_ready(FFs_14_io_d_rob_ready),
    .io_clear(FFs_14_io_clear)
  );
  prim_ff_cl_19 FFs_15 ( 
    .clock(FFs_15_clock),
    .reset(FFs_15_reset),
    .io_q_rob_type(FFs_15_io_q_rob_type),
    .io_q_rob_dest(FFs_15_io_q_rob_dest),
    .io_q_rob_value(FFs_15_io_q_rob_value),
    .io_q_rob_ready(FFs_15_io_q_rob_ready),
    .io_d_rob_type(FFs_15_io_d_rob_type),
    .io_d_rob_dest(FFs_15_io_d_rob_dest),
    .io_d_rob_value(FFs_15_io_d_rob_value),
    .io_d_rob_ready(FFs_15_io_d_rob_ready),
    .io_clear(FFs_15_io_clear)
  );
  assign io_enq_idx = h_ptr_io_q; 
  assign io_deq_data = {io_deq_data_hi,io_deq_data_lo}; 
  assign io_deq_idx = t_ptr_io_q; 
  assign io_empty = h_ptr_io_q == t_ptr_io_q; 
  assign io_full = _io_full_T_1 == t_ptr_io_q; 
  assign io_queue_data = {io_queue_data_hi,io_queue_data_lo}; 
  assign h_ptr_clock = clock;
  assign h_ptr_reset = reset;
  assign h_ptr_io_d = io_enq & ~io_full ? _io_full_T_1 : h_ptr_io_q; 
  assign h_ptr_io_clear = io_clear; 
  assign t_ptr_clock = clock;
  assign t_ptr_reset = reset;
  assign t_ptr_io_d = io_deq & ~io_empty ? _t_ptr_io_d_T_1 : t_ptr_io_q; 
  assign t_ptr_io_clear = io_clear; 
  assign FFs_0_clock = clock;
  assign FFs_0_reset = reset;
  assign FFs_0_io_d_rob_type = 4'h0 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_69; 
  assign FFs_0_io_d_rob_dest = 4'h0 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_68; 
  assign FFs_0_io_d_rob_value = 4'h0 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_67; 
  assign FFs_0_io_d_rob_ready = 4'h0 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_66; 
  assign FFs_0_io_clear = 4'h0 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_1_clock = clock;
  assign FFs_1_reset = reset;
  assign FFs_1_io_d_rob_type = 4'h1 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_78; 
  assign FFs_1_io_d_rob_dest = 4'h1 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_77; 
  assign FFs_1_io_d_rob_value = 4'h1 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_76; 
  assign FFs_1_io_d_rob_ready = 4'h1 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_75; 
  assign FFs_1_io_clear = 4'h1 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_2_clock = clock;
  assign FFs_2_reset = reset;
  assign FFs_2_io_d_rob_type = 4'h2 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_87; 
  assign FFs_2_io_d_rob_dest = 4'h2 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_86; 
  assign FFs_2_io_d_rob_value = 4'h2 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_85; 
  assign FFs_2_io_d_rob_ready = 4'h2 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_84; 
  assign FFs_2_io_clear = 4'h2 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_3_clock = clock;
  assign FFs_3_reset = reset;
  assign FFs_3_io_d_rob_type = 4'h3 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_96; 
  assign FFs_3_io_d_rob_dest = 4'h3 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_95; 
  assign FFs_3_io_d_rob_value = 4'h3 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_94; 
  assign FFs_3_io_d_rob_ready = 4'h3 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_93; 
  assign FFs_3_io_clear = 4'h3 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_4_clock = clock;
  assign FFs_4_reset = reset;
  assign FFs_4_io_d_rob_type = 4'h4 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_105; 
  assign FFs_4_io_d_rob_dest = 4'h4 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_104; 
  assign FFs_4_io_d_rob_value = 4'h4 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_103; 
  assign FFs_4_io_d_rob_ready = 4'h4 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_102; 
  assign FFs_4_io_clear = 4'h4 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_5_clock = clock;
  assign FFs_5_reset = reset;
  assign FFs_5_io_d_rob_type = 4'h5 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_114; 
  assign FFs_5_io_d_rob_dest = 4'h5 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_113; 
  assign FFs_5_io_d_rob_value = 4'h5 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_112; 
  assign FFs_5_io_d_rob_ready = 4'h5 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_111; 
  assign FFs_5_io_clear = 4'h5 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_6_clock = clock;
  assign FFs_6_reset = reset;
  assign FFs_6_io_d_rob_type = 4'h6 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_123; 
  assign FFs_6_io_d_rob_dest = 4'h6 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_122; 
  assign FFs_6_io_d_rob_value = 4'h6 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_121; 
  assign FFs_6_io_d_rob_ready = 4'h6 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_120; 
  assign FFs_6_io_clear = 4'h6 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_7_clock = clock;
  assign FFs_7_reset = reset;
  assign FFs_7_io_d_rob_type = 4'h7 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_132; 
  assign FFs_7_io_d_rob_dest = 4'h7 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_131; 
  assign FFs_7_io_d_rob_value = 4'h7 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_130; 
  assign FFs_7_io_d_rob_ready = 4'h7 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_129; 
  assign FFs_7_io_clear = 4'h7 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_8_clock = clock;
  assign FFs_8_reset = reset;
  assign FFs_8_io_d_rob_type = 4'h8 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_141; 
  assign FFs_8_io_d_rob_dest = 4'h8 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_140; 
  assign FFs_8_io_d_rob_value = 4'h8 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_139; 
  assign FFs_8_io_d_rob_ready = 4'h8 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_138; 
  assign FFs_8_io_clear = 4'h8 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_9_clock = clock;
  assign FFs_9_reset = reset;
  assign FFs_9_io_d_rob_type = 4'h9 == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_150; 
  assign FFs_9_io_d_rob_dest = 4'h9 == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_149; 
  assign FFs_9_io_d_rob_value = 4'h9 == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_148; 
  assign FFs_9_io_d_rob_ready = 4'h9 == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_147; 
  assign FFs_9_io_clear = 4'h9 == io_deq_idx & _T_4 | io_clear; 
  assign FFs_10_clock = clock;
  assign FFs_10_reset = reset;
  assign FFs_10_io_d_rob_type = 4'ha == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_159; 
  assign FFs_10_io_d_rob_dest = 4'ha == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_158; 
  assign FFs_10_io_d_rob_value = 4'ha == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_157; 
  assign FFs_10_io_d_rob_ready = 4'ha == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_156; 
  assign FFs_10_io_clear = 4'ha == io_deq_idx & _T_4 | io_clear; 
  assign FFs_11_clock = clock;
  assign FFs_11_reset = reset;
  assign FFs_11_io_d_rob_type = 4'hb == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_168; 
  assign FFs_11_io_d_rob_dest = 4'hb == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_167; 
  assign FFs_11_io_d_rob_value = 4'hb == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_166; 
  assign FFs_11_io_d_rob_ready = 4'hb == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_165; 
  assign FFs_11_io_clear = 4'hb == io_deq_idx & _T_4 | io_clear; 
  assign FFs_12_clock = clock;
  assign FFs_12_reset = reset;
  assign FFs_12_io_d_rob_type = 4'hc == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_177; 
  assign FFs_12_io_d_rob_dest = 4'hc == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_176; 
  assign FFs_12_io_d_rob_value = 4'hc == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_175; 
  assign FFs_12_io_d_rob_ready = 4'hc == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_174; 
  assign FFs_12_io_clear = 4'hc == io_deq_idx & _T_4 | io_clear; 
  assign FFs_13_clock = clock;
  assign FFs_13_reset = reset;
  assign FFs_13_io_d_rob_type = 4'hd == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_186; 
  assign FFs_13_io_d_rob_dest = 4'hd == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_185; 
  assign FFs_13_io_d_rob_value = 4'hd == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_184; 
  assign FFs_13_io_d_rob_ready = 4'hd == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_183; 
  assign FFs_13_io_clear = 4'hd == io_deq_idx & _T_4 | io_clear; 
  assign FFs_14_clock = clock;
  assign FFs_14_reset = reset;
  assign FFs_14_io_d_rob_type = 4'he == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_195; 
  assign FFs_14_io_d_rob_dest = 4'he == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_194; 
  assign FFs_14_io_d_rob_value = 4'he == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_193; 
  assign FFs_14_io_d_rob_ready = 4'he == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_192; 
  assign FFs_14_io_clear = 4'he == io_deq_idx & _T_4 | io_clear; 
  assign FFs_15_clock = clock;
  assign FFs_15_reset = reset;
  assign FFs_15_io_d_rob_type = 4'hf == io_enq_idx & _T_1 ? io_enq_data[66:65] : _GEN_204; 
  assign FFs_15_io_d_rob_dest = 4'hf == io_enq_idx & _T_1 ? io_enq_data[64:33] : _GEN_203; 
  assign FFs_15_io_d_rob_value = 4'hf == io_enq_idx & _T_1 ? io_enq_data[32:1] : _GEN_202; 
  assign FFs_15_io_d_rob_ready = 4'hf == io_enq_idx & _T_1 ? io_enq_data[0] : _GEN_201; 
  assign FFs_15_io_clear = 4'hf == io_deq_idx & _T_4 | io_clear; 
endmodule
module FIFO_ROB(
  input           clock,
  input           reset,
  input           io_clear, 
  input           io_enq, 
  input  [66:0]   io_enq_data, 
  input           io_deq, 
  output [66:0]   io_deq_data, 
  output          io_empty, 
  output          io_full, 
  output [4:0]    io_enq_idx, 
  output [4:0]    io_deq_idx, 
  output [1138:0] io_queue_data, 
  input  [16:0]   io_update_entry, 
  input  [1138:0] io_update_entry_data 
);
  wire  mFIFO_clock; 
  wire  mFIFO_reset; 
  wire  mFIFO_io_clear; 
  wire  mFIFO_io_enq; 
  wire [66:0] mFIFO_io_enq_data; 
  wire [3:0] mFIFO_io_enq_idx; 
  wire  mFIFO_io_deq; 
  wire [66:0] mFIFO_io_deq_data; 
  wire [3:0] mFIFO_io_deq_idx; 
  wire  mFIFO_io_empty; 
  wire  mFIFO_io_full; 
  wire [1071:0] mFIFO_io_queue_data; 
  wire [15:0] mFIFO_io_update_entry; 
  wire [1071:0] mFIFO_io_update_entry_data; 
  FIFO_2 mFIFO ( 
    .clock(mFIFO_clock),
    .reset(mFIFO_reset),
    .io_clear(mFIFO_io_clear),
    .io_enq(mFIFO_io_enq),
    .io_enq_data(mFIFO_io_enq_data),
    .io_enq_idx(mFIFO_io_enq_idx),
    .io_deq(mFIFO_io_deq),
    .io_deq_data(mFIFO_io_deq_data),
    .io_deq_idx(mFIFO_io_deq_idx),
    .io_empty(mFIFO_io_empty),
    .io_full(mFIFO_io_full),
    .io_queue_data(mFIFO_io_queue_data),
    .io_update_entry(mFIFO_io_update_entry),
    .io_update_entry_data(mFIFO_io_update_entry_data)
  );
  assign io_deq_data = mFIFO_io_deq_data; 
  assign io_empty = mFIFO_io_empty; 
  assign io_full = mFIFO_io_full; 
  assign io_enq_idx = mFIFO_io_enq_idx + 4'h1; 
  assign io_deq_idx = mFIFO_io_deq_idx + 4'h1; 
  assign io_queue_data = {mFIFO_io_queue_data,67'h0}; 
  assign mFIFO_clock = clock;
  assign mFIFO_reset = reset;
  assign mFIFO_io_clear = io_clear; 
  assign mFIFO_io_enq = io_enq; 
  assign mFIFO_io_enq_data = io_enq_data; 
  assign mFIFO_io_deq = io_deq; 
  assign mFIFO_io_update_entry = io_update_entry[16:1]; 
  assign mFIFO_io_update_entry_data = io_update_entry_data[1138:67]; 
endmodule
module prim_ff_cl_36(
  input         clock,
  input         reset,
  output        io_q_valid, 
  output [31:0] io_q_result, 
  output [4:0]  io_q_dest, 
  input         io_d_valid, 
  input  [31:0] io_d_result, 
  input  [4:0]  io_d_dest, 
  input         io_clear 
);
  reg  m_reg_valid; 
  reg [31:0] m_reg_result; 
  reg [4:0] m_reg_dest; 
  assign io_q_valid = m_reg_valid; 
  assign io_q_result = m_reg_result; 
  assign io_q_dest = m_reg_dest; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_valid <= 1'h0; 
    end else if (io_clear) begin 
      m_reg_valid <= 1'h0;
    end else begin
      m_reg_valid <= io_d_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_result <= 32'h0; 
    end else if (io_clear) begin 
      m_reg_result <= 32'h0;
    end else begin
      m_reg_result <= io_d_result;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_dest <= 5'h0; 
    end else if (io_clear) begin 
      m_reg_dest <= 5'h0;
    end else begin
      m_reg_dest <= io_d_dest;
    end
  end
endmodule
module CDB(
  input         clock,
  input         reset,
  input         io_clear, 
  input         io_int_valid, 
  output        io_int_ready, 
  input  [31:0] io_int_result, 
  input  [4:0]  io_int_dest, 
  input         io_muldiv_valid, 
  output        io_muldiv_ready, 
  input  [31:0] io_muldiv_result, 
  input  [4:0]  io_muldiv_dest, 
  input         io_mem_valid, 
  output        io_mem_ready, 
  input  [31:0] io_mem_result, 
  input  [4:0]  io_mem_dest, 
  output        io_cdb_valid, 
  output [31:0] io_cdb_result, 
  output [4:0]  io_cdb_dest 
);
  wire  mState_clock; 
  wire  mState_reset; 
  wire [1:0] mState_io_q; 
  wire [1:0] mState_io_d; 
  wire  mState_io_clear; 
  wire  out_clock; 
  wire  out_reset; 
  wire  out_io_q_valid; 
  wire [31:0] out_io_q_result; 
  wire [4:0] out_io_q_dest; 
  wire  out_io_d_valid; 
  wire [31:0] out_io_d_result; 
  wire [4:0] out_io_d_dest; 
  wire  out_io_clear; 
  wire  m_mem_rcy_clock; 
  wire  m_mem_rcy_reset; 
  wire  m_mem_rcy_io_q_valid; 
  wire [31:0] m_mem_rcy_io_q_result; 
  wire [4:0] m_mem_rcy_io_q_dest; 
  wire  m_mem_rcy_io_d_valid; 
  wire [31:0] m_mem_rcy_io_d_result; 
  wire [4:0] m_mem_rcy_io_d_dest; 
  wire  m_mem_rcy_io_clear; 
  wire  m_int_rcy_clock; 
  wire  m_int_rcy_reset; 
  wire  m_int_rcy_io_q_valid; 
  wire [31:0] m_int_rcy_io_q_result; 
  wire [4:0] m_int_rcy_io_q_dest; 
  wire  m_int_rcy_io_d_valid; 
  wire [31:0] m_int_rcy_io_d_result; 
  wire [4:0] m_int_rcy_io_d_dest; 
  wire  m_int_rcy_io_clear; 
  wire  _io_muldiv_ready_T_2 = mState_io_q == 2'h0; 
  wire  _io_mem_ready_T = ~io_muldiv_valid; 
  wire  _io_int_ready_T_7 = io_int_valid & ~io_mem_valid & _io_mem_ready_T & _io_muldiv_ready_T_2; 
  wire [1:0] mStateEnum = mState_io_q; 
  wire [4:0] _GEN_0 = io_int_valid ? io_int_dest : out_io_q_dest; 
  wire [31:0] _GEN_1 = io_int_valid ? io_int_result : out_io_q_result; 
  wire [4:0] _GEN_3 = io_mem_valid ? io_mem_dest : _GEN_0; 
  wire [31:0] _GEN_4 = io_mem_valid ? io_mem_result : _GEN_1; 
  wire  _GEN_5 = io_mem_valid | io_int_valid; 
  wire [4:0] _GEN_7 = io_muldiv_valid ? io_muldiv_dest : _GEN_3; 
  wire [31:0] _GEN_8 = io_muldiv_valid ? io_muldiv_result : _GEN_4; 
  wire  _GEN_9 = io_muldiv_valid | _GEN_5; 
  wire  _T_10 = io_muldiv_valid & io_mem_valid; 
  wire  _T_13 = io_int_valid & (io_mem_valid | io_muldiv_valid); 
  wire [1:0] _GEN_11 = io_int_valid & (io_mem_valid | io_muldiv_valid) ? 2'h2 : 2'h0; 
  wire [4:0] _GEN_12 = io_int_valid & (io_mem_valid | io_muldiv_valid) ? io_int_dest : m_int_rcy_io_q_dest; 
  wire [31:0] _GEN_13 = io_int_valid & (io_mem_valid | io_muldiv_valid) ? io_int_result : m_int_rcy_io_q_result; 
  wire [1:0] _GEN_15 = io_muldiv_valid & io_mem_valid ? 2'h1 : _GEN_11; 
  wire [4:0] _GEN_16 = io_muldiv_valid & io_mem_valid ? io_mem_dest : m_mem_rcy_io_q_dest; 
  wire [31:0] _GEN_17 = io_muldiv_valid & io_mem_valid ? io_mem_result : m_mem_rcy_io_q_result; 
  wire [4:0] _GEN_19 = io_muldiv_valid & io_mem_valid ? m_int_rcy_io_q_dest : _GEN_12; 
  wire [31:0] _GEN_20 = io_muldiv_valid & io_mem_valid ? m_int_rcy_io_q_result : _GEN_13; 
  wire  _GEN_21 = io_muldiv_valid & io_mem_valid ? 1'h0 : _T_13; 
  wire [1:0] _GEN_22 = m_int_rcy_io_q_valid ? 2'h2 : 2'h0; 
  wire [4:0] _GEN_23 = 2'h2 == mStateEnum ? m_int_rcy_io_q_dest : out_io_q_dest; 
  wire [31:0] _GEN_24 = 2'h2 == mStateEnum ? m_int_rcy_io_q_result : out_io_q_result; 
  wire [1:0] _GEN_26 = 2'h2 == mStateEnum ? 2'h0 : mState_io_q; 
  wire [4:0] _GEN_27 = 2'h1 == mStateEnum ? m_mem_rcy_io_q_dest : _GEN_23; 
  wire [31:0] _GEN_28 = 2'h1 == mStateEnum ? m_mem_rcy_io_q_result : _GEN_24; 
  wire  _GEN_29 = 2'h1 == mStateEnum | 2'h2 == mStateEnum; 
  wire [1:0] _GEN_31 = 2'h1 == mStateEnum ? _GEN_22 : _GEN_26; 
  prim_ff_cl_5 mState ( 
    .clock(mState_clock),
    .reset(mState_reset),
    .io_q(mState_io_q),
    .io_d(mState_io_d),
    .io_clear(mState_io_clear)
  );
  prim_ff_cl_36 out ( 
    .clock(out_clock),
    .reset(out_reset),
    .io_q_valid(out_io_q_valid),
    .io_q_result(out_io_q_result),
    .io_q_dest(out_io_q_dest),
    .io_d_valid(out_io_d_valid),
    .io_d_result(out_io_d_result),
    .io_d_dest(out_io_d_dest),
    .io_clear(out_io_clear)
  );
  prim_ff_cl_36 m_mem_rcy ( 
    .clock(m_mem_rcy_clock),
    .reset(m_mem_rcy_reset),
    .io_q_valid(m_mem_rcy_io_q_valid),
    .io_q_result(m_mem_rcy_io_q_result),
    .io_q_dest(m_mem_rcy_io_q_dest),
    .io_d_valid(m_mem_rcy_io_d_valid),
    .io_d_result(m_mem_rcy_io_d_result),
    .io_d_dest(m_mem_rcy_io_d_dest),
    .io_clear(m_mem_rcy_io_clear)
  );
  prim_ff_cl_36 m_int_rcy ( 
    .clock(m_int_rcy_clock),
    .reset(m_int_rcy_reset),
    .io_q_valid(m_int_rcy_io_q_valid),
    .io_q_result(m_int_rcy_io_q_result),
    .io_q_dest(m_int_rcy_io_q_dest),
    .io_d_valid(m_int_rcy_io_d_valid),
    .io_d_result(m_int_rcy_io_d_result),
    .io_d_dest(m_int_rcy_io_d_dest),
    .io_clear(m_int_rcy_io_clear)
  );
  assign io_int_ready = _io_int_ready_T_7 | mState_io_q == 2'h2; 
  assign io_muldiv_ready = io_muldiv_valid & mState_io_q == 2'h0; 
  assign io_mem_ready = io_mem_valid & ~io_muldiv_valid & _io_muldiv_ready_T_2 | mState_io_q == 2'h1; 
  assign io_cdb_valid = out_io_q_valid; 
  assign io_cdb_result = out_io_q_result; 
  assign io_cdb_dest = out_io_q_dest; 
  assign mState_clock = clock;
  assign mState_reset = reset;
  assign mState_io_d = 2'h0 == mStateEnum ? _GEN_15 : _GEN_31; 
  assign mState_io_clear = io_clear; 
  assign out_clock = clock;
  assign out_reset = reset;
  assign out_io_d_valid = 2'h0 == mStateEnum ? _GEN_9 : _GEN_29; 
  assign out_io_d_result = 2'h0 == mStateEnum ? _GEN_8 : _GEN_28; 
  assign out_io_d_dest = 2'h0 == mStateEnum ? _GEN_7 : _GEN_27; 
  assign out_io_clear = io_clear; 
  assign m_mem_rcy_clock = clock;
  assign m_mem_rcy_reset = reset;
  assign m_mem_rcy_io_d_valid = 2'h0 == mStateEnum & _T_10; 
  assign m_mem_rcy_io_d_result = 2'h0 == mStateEnum ? _GEN_17 : m_mem_rcy_io_q_result; 
  assign m_mem_rcy_io_d_dest = 2'h0 == mStateEnum ? _GEN_16 : m_mem_rcy_io_q_dest; 
  assign m_mem_rcy_io_clear = io_clear; 
  assign m_int_rcy_clock = clock;
  assign m_int_rcy_reset = reset;
  assign m_int_rcy_io_d_valid = 2'h0 == mStateEnum & _GEN_21; 
  assign m_int_rcy_io_d_result = 2'h0 == mStateEnum ? _GEN_20 : m_int_rcy_io_q_result; 
  assign m_int_rcy_io_d_dest = 2'h0 == mStateEnum ? _GEN_19 : m_int_rcy_io_q_dest; 
  assign m_int_rcy_io_clear = io_clear; 
endmodule
module IntOp(
  input         clock,
  input         reset,
  input         io_clear, 
  input         io_in_valid, 
  input  [31:0] io_in_in1, 
  input  [31:0] io_in_in2, 
  input         io_in_op_store, 
  input         io_in_op_load, 
  input         io_in_op_muldivb_s, 
  input         io_in_op_muldiva_s, 
  input         io_in_op_div, 
  input         io_in_op_mul, 
  input         io_in_op_equal, 
  input         io_in_op_large, 
  input         io_in_op_less, 
  input         io_in_op_jr, 
  input         io_in_op_br, 
  input         io_in_op_sra, 
  input         io_in_op_srl, 
  input         io_in_op_sll, 
  input         io_in_op_sub, 
  input         io_in_op_add, 
  input         io_in_op_set, 
  input         io_in_op_xor, 
  input         io_in_op_or, 
  input         io_in_op_and, 
  input  [4:0]  io_in_dest, 
  output        io_out_valid, 
  output [31:0] io_out_result, 
  output [4:0]  io_out_dest 
);
  wire  uOp_clock; 
  wire  uOp_reset; 
  wire  uOp_clear; 
  wire  uOp_valid; 
  wire [19:0] uOp_op; 
  wire [31:0] uOp_in_1; 
  wire [31:0] uOp_in_2; 
  wire [4:0] uOp_RS_idx_i; 
  wire  uOp_result_valid; 
  wire [31:0] uOp_result; 
  wire [4:0] uOp_RS_idx_o; 
  wire  uOp_branch_finish; 
  wire  uOp_branch_true; 
  wire [9:0] uOp_io_op_lo = {io_in_op_br,io_in_op_sra,io_in_op_srl,io_in_op_sll,io_in_op_sub,io_in_op_add,io_in_op_set,
    io_in_op_xor,io_in_op_or,io_in_op_and}; 
  wire [9:0] uOp_io_op_hi = {io_in_op_store,io_in_op_load,io_in_op_muldivb_s,io_in_op_muldiva_s,io_in_op_div,
    io_in_op_mul,io_in_op_equal,io_in_op_large,io_in_op_less,io_in_op_jr}; 
  integer_operation uOp ( 
    .clock(uOp_clock),
    .reset(uOp_reset),
    .clear(uOp_clear),
    .valid(uOp_valid),
    .op(uOp_op),
    .in_1(uOp_in_1),
    .in_2(uOp_in_2),
    .RS_idx_i(uOp_RS_idx_i),
    .result_valid(uOp_result_valid),
    .result(uOp_result),
    .RS_idx_o(uOp_RS_idx_o),
    .branch_finish(uOp_branch_finish),
    .branch_true(uOp_branch_true)
  );
  assign io_out_valid = uOp_result_valid; 
  assign io_out_result = uOp_result; 
  assign io_out_dest = uOp_RS_idx_o; 
  assign uOp_clock = clock; 
  assign uOp_reset = reset; 
  assign uOp_clear = io_clear; 
  assign uOp_valid = io_in_valid; 
  assign uOp_op = {uOp_io_op_hi,uOp_io_op_lo}; 
  assign uOp_in_1 = io_in_in1; 
  assign uOp_in_2 = io_in_in2; 
  assign uOp_RS_idx_i = io_in_dest; 
endmodule
module MulDivOp(
  input         clock,
  input         reset,
  input         io_clear, 
  input         io_in_valid, 
  input  [31:0] io_in_in1, 
  input  [31:0] io_in_in2, 
  input         io_in_op_muldivb_s, 
  input         io_in_op_muldiva_s, 
  input         io_in_op_mul, 
  input  [4:0]  io_in_dest, 
  output        io_out_valid, 
  output [31:0] io_out_result, 
  output [4:0]  io_out_dest 
);
  wire  uOp_clock; 
  wire  uOp_reset; 
  wire  uOp_clear; 
  wire  uOp_valid; 
  wire  uOp_mul1_div0; 
  wire [1:0] uOp_in_sign; 
  wire [31:0] uOp_operation_in_1; 
  wire [31:0] uOp_operation_in_2; 
  wire [4:0] uOp_RS_idx_i; 
  wire  uOp_result_valid; 
  wire [31:0] uOp_result; 
  wire [4:0] uOp_RS_idx_o; 
  muldiv_operation #(.DIV_CYCLE(10), .MUL_CYCLE(6)) uOp ( 
    .clock(uOp_clock),
    .reset(uOp_reset),
    .clear(uOp_clear),
    .valid(uOp_valid),
    .mul1_div0(uOp_mul1_div0),
    .in_sign(uOp_in_sign),
    .operation_in_1(uOp_operation_in_1),
    .operation_in_2(uOp_operation_in_2),
    .RS_idx_i(uOp_RS_idx_i),
    .result_valid(uOp_result_valid),
    .result(uOp_result),
    .RS_idx_o(uOp_RS_idx_o)
  );
  assign io_out_valid = uOp_result_valid; 
  assign io_out_result = uOp_result; 
  assign io_out_dest = uOp_RS_idx_o; 
  assign uOp_clock = clock; 
  assign uOp_reset = reset; 
  assign uOp_clear = io_clear; 
  assign uOp_valid = io_in_valid; 
  assign uOp_mul1_div0 = io_in_op_mul; 
  assign uOp_in_sign = {io_in_op_muldivb_s,io_in_op_muldiva_s}; 
  assign uOp_operation_in_1 = io_in_in1; 
  assign uOp_operation_in_2 = io_in_in2; 
  assign uOp_RS_idx_i = io_in_dest; 
endmodule
module prim_ff_cl_39(
  input         clock,
  input         reset,
  output [31:0] io_q, 
  input  [31:0] io_d, 
  input         io_clear 
);
  reg [31:0] m_reg; 
  assign io_q = m_reg; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg <= 32'h0; 
    end else if (io_clear) begin 
      m_reg <= 32'h0;
    end else begin
      m_reg <= io_d;
    end
  end
endmodule
module prim_ff_cl_71(
  input        clock,
  input        reset,
  output       io_q_busy, 
  output [4:0] io_q_reorder, 
  input        io_d_busy, 
  input  [4:0] io_d_reorder, 
  input        io_clear 
);
  reg  m_reg_busy; 
  reg [4:0] m_reg_reorder; 
  assign io_q_busy = m_reg_busy; 
  assign io_q_reorder = m_reg_reorder; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_busy <= 1'h0; 
    end else if (io_clear) begin 
      m_reg_busy <= 1'h0;
    end else begin
      m_reg_busy <= io_d_busy;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg_reorder <= 5'h0; 
    end else if (io_clear) begin 
      m_reg_reorder <= 5'h0;
    end else begin
      m_reg_reorder <= io_d_reorder;
    end
  end
endmodule
module prim_ff_cl_103(
  input   clock,
  input   reset,
  output  io_q, 
  input   io_d, 
  input   io_clear 
);
  reg  m_reg; 
  assign io_q = m_reg; 
  always @(posedge clock or posedge reset) begin
    if (reset) begin 
      m_reg <= 1'h0; 
    end else if (io_clear) begin 
      m_reg <= 1'h0;
    end else begin
      m_reg <= io_d;
    end
  end
endmodule
module RiscvCoreTop(
  input         clock,
  input         reset,
  input         decoder_if_inst_valid, 
  input         decoder_if_exe_op_store, 
  input         decoder_if_exe_op_load, 
  input         decoder_if_exe_op_muldivb_s, 
  input         decoder_if_exe_op_muldiva_s, 
  input         decoder_if_exe_op_div, 
  input         decoder_if_exe_op_mul, 
  input         decoder_if_exe_op_equal, 
  input         decoder_if_exe_op_large, 
  input         decoder_if_exe_op_less, 
  input         decoder_if_exe_op_jr, 
  input         decoder_if_exe_op_br, 
  input         decoder_if_exe_op_sra, 
  input         decoder_if_exe_op_srl, 
  input         decoder_if_exe_op_sll, 
  input         decoder_if_exe_op_sub, 
  input         decoder_if_exe_op_add, 
  input         decoder_if_exe_op_set, 
  input         decoder_if_exe_op_xor, 
  input         decoder_if_exe_op_or, 
  input         decoder_if_exe_op_and, 
  input  [31:0] decoder_if_imm, 
  input         decoder_if_imm_valid, 
  input  [31:0] decoder_if_pc_out, 
  input         decoder_if_pc_valid, 
  input  [4:0]  decoder_if_rs_idx, 
  input         decoder_if_rs_idx_valid, 
  input  [4:0]  decoder_if_rt_idx, 
  input         decoder_if_rt_idx_valid, 
  input  [4:0]  decoder_if_rd_idx, 
  input         decoder_if_rd_idx_valid, 
  output        fetcher_if_stall_fetch, 
  output        fetcher_if_re_jump_en, 
  output [31:0] fetcher_if_re_jump_addr, 
  output [4:0]  datamem_if_RS_idx_i, 
  input  [4:0]  datamem_if_RS_idx_o, 
  output        datamem_if_st_valid, 
  input         datamem_if_st_ready, 
  output [31:0] datamem_if_st_addr, 
  output [31:0] datamem_if_st_data, 
  output        datamem_if_ld_valid, 
  input         datamem_if_ld_ready, 
  output [31:0] datamem_if_ld_addr, 
  input  [31:0] datamem_if_ld_data, 
  input         datamem_if_ld_data_valid 
);
  wire  uIntergerRS__clock; 
  wire  uIntergerRS__reset; 
  wire  uIntergerRS__io_clear; 
  wire  uIntergerRS__io_enq; 
  wire [131:0] uIntergerRS__io_enq_data; 
  wire  uIntergerRS__io_deq; 
  wire [3:0] uIntergerRS__io_deq_cond; 
  wire [131:0] uIntergerRS__io_deq_data; 
  wire  uIntergerRS__io_empty; 
  wire  uIntergerRS__io_full; 
  wire [527:0] uIntergerRS__io_queue_data; 
  wire [3:0] uIntergerRS__io_update_entry; 
  wire [527:0] uIntergerRS__io_update_entry_data; 
  wire  uMulDivRS__clock; 
  wire  uMulDivRS__reset; 
  wire  uMulDivRS__io_clear; 
  wire  uMulDivRS__io_enq; 
  wire [131:0] uMulDivRS__io_enq_data; 
  wire [1:0] uMulDivRS__io_enq_idx; 
  wire  uMulDivRS__io_deq; 
  wire [131:0] uMulDivRS__io_deq_data; 
  wire [1:0] uMulDivRS__io_deq_idx; 
  wire  uMulDivRS__io_empty; 
  wire  uMulDivRS__io_full; 
  wire [527:0] uMulDivRS__io_queue_data; 
  wire [3:0] uMulDivRS__io_update_entry; 
  wire [527:0] uMulDivRS__io_update_entry_data; 
  wire  uLoadStoreRS__clock; 
  wire  uLoadStoreRS__reset; 
  wire  uLoadStoreRS__io_clear; 
  wire  uLoadStoreRS__io_enq; 
  wire [131:0] uLoadStoreRS__io_enq_data; 
  wire [1:0] uLoadStoreRS__io_enq_idx; 
  wire  uLoadStoreRS__io_deq; 
  wire [131:0] uLoadStoreRS__io_deq_data; 
  wire [1:0] uLoadStoreRS__io_deq_idx; 
  wire  uLoadStoreRS__io_empty; 
  wire  uLoadStoreRS__io_full; 
  wire [527:0] uLoadStoreRS__io_queue_data; 
  wire [3:0] uLoadStoreRS__io_update_entry; 
  wire [527:0] uLoadStoreRS__io_update_entry_data; 
  wire  uROB__clock; 
  wire  uROB__reset; 
  wire  uROB__io_clear; 
  wire  uROB__io_enq; 
  wire [66:0] uROB__io_enq_data; 
  wire  uROB__io_deq; 
  wire [66:0] uROB__io_deq_data; 
  wire  uROB__io_empty; 
  wire  uROB__io_full; 
  wire [4:0] uROB__io_enq_idx; 
  wire [4:0] uROB__io_deq_idx; 
  wire [1138:0] uROB__io_queue_data; 
  wire [16:0] uROB__io_update_entry; 
  wire [1138:0] uROB__io_update_entry_data; 
  wire  uCDB_clock; 
  wire  uCDB_reset; 
  wire  uCDB_io_clear; 
  wire  uCDB_io_int_valid; 
  wire  uCDB_io_int_ready; 
  wire [31:0] uCDB_io_int_result; 
  wire [4:0] uCDB_io_int_dest; 
  wire  uCDB_io_muldiv_valid; 
  wire  uCDB_io_muldiv_ready; 
  wire [31:0] uCDB_io_muldiv_result; 
  wire [4:0] uCDB_io_muldiv_dest; 
  wire  uCDB_io_mem_valid; 
  wire  uCDB_io_mem_ready; 
  wire [31:0] uCDB_io_mem_result; 
  wire [4:0] uCDB_io_mem_dest; 
  wire  uCDB_io_cdb_valid; 
  wire [31:0] uCDB_io_cdb_result; 
  wire [4:0] uCDB_io_cdb_dest; 
  wire  uIntOp_clock; 
  wire  uIntOp_reset; 
  wire  uIntOp_io_clear; 
  wire  uIntOp_io_in_valid; 
  wire [31:0] uIntOp_io_in_in1; 
  wire [31:0] uIntOp_io_in_in2; 
  wire  uIntOp_io_in_op_store; 
  wire  uIntOp_io_in_op_load; 
  wire  uIntOp_io_in_op_muldivb_s; 
  wire  uIntOp_io_in_op_muldiva_s; 
  wire  uIntOp_io_in_op_div; 
  wire  uIntOp_io_in_op_mul; 
  wire  uIntOp_io_in_op_equal; 
  wire  uIntOp_io_in_op_large; 
  wire  uIntOp_io_in_op_less; 
  wire  uIntOp_io_in_op_jr; 
  wire  uIntOp_io_in_op_br; 
  wire  uIntOp_io_in_op_sra; 
  wire  uIntOp_io_in_op_srl; 
  wire  uIntOp_io_in_op_sll; 
  wire  uIntOp_io_in_op_sub; 
  wire  uIntOp_io_in_op_add; 
  wire  uIntOp_io_in_op_set; 
  wire  uIntOp_io_in_op_xor; 
  wire  uIntOp_io_in_op_or; 
  wire  uIntOp_io_in_op_and; 
  wire [4:0] uIntOp_io_in_dest; 
  wire  uIntOp_io_out_valid; 
  wire [31:0] uIntOp_io_out_result; 
  wire [4:0] uIntOp_io_out_dest; 
  wire  uMulDivOp_clock; 
  wire  uMulDivOp_reset; 
  wire  uMulDivOp_io_clear; 
  wire  uMulDivOp_io_in_valid; 
  wire [31:0] uMulDivOp_io_in_in1; 
  wire [31:0] uMulDivOp_io_in_in2; 
  wire  uMulDivOp_io_in_op_muldivb_s; 
  wire  uMulDivOp_io_in_op_muldiva_s; 
  wire  uMulDivOp_io_in_op_mul; 
  wire [4:0] uMulDivOp_io_in_dest; 
  wire  uMulDivOp_io_out_valid; 
  wire [31:0] uMulDivOp_io_out_result; 
  wire [4:0] uMulDivOp_io_out_dest; 
  wire  uRegFile_0_clock; 
  wire  uRegFile_0_reset; 
  wire [31:0] uRegFile_0_io_q; 
  wire [31:0] uRegFile_0_io_d; 
  wire  uRegFile_0_io_clear; 
  wire  uRegFile_1_clock; 
  wire  uRegFile_1_reset; 
  wire [31:0] uRegFile_1_io_q; 
  wire [31:0] uRegFile_1_io_d; 
  wire  uRegFile_1_io_clear; 
  wire  uRegFile_2_clock; 
  wire  uRegFile_2_reset; 
  wire [31:0] uRegFile_2_io_q; 
  wire [31:0] uRegFile_2_io_d; 
  wire  uRegFile_2_io_clear; 
  wire  uRegFile_3_clock; 
  wire  uRegFile_3_reset; 
  wire [31:0] uRegFile_3_io_q; 
  wire [31:0] uRegFile_3_io_d; 
  wire  uRegFile_3_io_clear; 
  wire  uRegFile_4_clock; 
  wire  uRegFile_4_reset; 
  wire [31:0] uRegFile_4_io_q; 
  wire [31:0] uRegFile_4_io_d; 
  wire  uRegFile_4_io_clear; 
  wire  uRegFile_5_clock; 
  wire  uRegFile_5_reset; 
  wire [31:0] uRegFile_5_io_q; 
  wire [31:0] uRegFile_5_io_d; 
  wire  uRegFile_5_io_clear; 
  wire  uRegFile_6_clock; 
  wire  uRegFile_6_reset; 
  wire [31:0] uRegFile_6_io_q; 
  wire [31:0] uRegFile_6_io_d; 
  wire  uRegFile_6_io_clear; 
  wire  uRegFile_7_clock; 
  wire  uRegFile_7_reset; 
  wire [31:0] uRegFile_7_io_q; 
  wire [31:0] uRegFile_7_io_d; 
  wire  uRegFile_7_io_clear; 
  wire  uRegFile_8_clock; 
  wire  uRegFile_8_reset; 
  wire [31:0] uRegFile_8_io_q; 
  wire [31:0] uRegFile_8_io_d; 
  wire  uRegFile_8_io_clear; 
  wire  uRegFile_9_clock; 
  wire  uRegFile_9_reset; 
  wire [31:0] uRegFile_9_io_q; 
  wire [31:0] uRegFile_9_io_d; 
  wire  uRegFile_9_io_clear; 
  wire  uRegFile_10_clock; 
  wire  uRegFile_10_reset; 
  wire [31:0] uRegFile_10_io_q; 
  wire [31:0] uRegFile_10_io_d; 
  wire  uRegFile_10_io_clear; 
  wire  uRegFile_11_clock; 
  wire  uRegFile_11_reset; 
  wire [31:0] uRegFile_11_io_q; 
  wire [31:0] uRegFile_11_io_d; 
  wire  uRegFile_11_io_clear; 
  wire  uRegFile_12_clock; 
  wire  uRegFile_12_reset; 
  wire [31:0] uRegFile_12_io_q; 
  wire [31:0] uRegFile_12_io_d; 
  wire  uRegFile_12_io_clear; 
  wire  uRegFile_13_clock; 
  wire  uRegFile_13_reset; 
  wire [31:0] uRegFile_13_io_q; 
  wire [31:0] uRegFile_13_io_d; 
  wire  uRegFile_13_io_clear; 
  wire  uRegFile_14_clock; 
  wire  uRegFile_14_reset; 
  wire [31:0] uRegFile_14_io_q; 
  wire [31:0] uRegFile_14_io_d; 
  wire  uRegFile_14_io_clear; 
  wire  uRegFile_15_clock; 
  wire  uRegFile_15_reset; 
  wire [31:0] uRegFile_15_io_q; 
  wire [31:0] uRegFile_15_io_d; 
  wire  uRegFile_15_io_clear; 
  wire  uRegFile_16_clock; 
  wire  uRegFile_16_reset; 
  wire [31:0] uRegFile_16_io_q; 
  wire [31:0] uRegFile_16_io_d; 
  wire  uRegFile_16_io_clear; 
  wire  uRegFile_17_clock; 
  wire  uRegFile_17_reset; 
  wire [31:0] uRegFile_17_io_q; 
  wire [31:0] uRegFile_17_io_d; 
  wire  uRegFile_17_io_clear; 
  wire  uRegFile_18_clock; 
  wire  uRegFile_18_reset; 
  wire [31:0] uRegFile_18_io_q; 
  wire [31:0] uRegFile_18_io_d; 
  wire  uRegFile_18_io_clear; 
  wire  uRegFile_19_clock; 
  wire  uRegFile_19_reset; 
  wire [31:0] uRegFile_19_io_q; 
  wire [31:0] uRegFile_19_io_d; 
  wire  uRegFile_19_io_clear; 
  wire  uRegFile_20_clock; 
  wire  uRegFile_20_reset; 
  wire [31:0] uRegFile_20_io_q; 
  wire [31:0] uRegFile_20_io_d; 
  wire  uRegFile_20_io_clear; 
  wire  uRegFile_21_clock; 
  wire  uRegFile_21_reset; 
  wire [31:0] uRegFile_21_io_q; 
  wire [31:0] uRegFile_21_io_d; 
  wire  uRegFile_21_io_clear; 
  wire  uRegFile_22_clock; 
  wire  uRegFile_22_reset; 
  wire [31:0] uRegFile_22_io_q; 
  wire [31:0] uRegFile_22_io_d; 
  wire  uRegFile_22_io_clear; 
  wire  uRegFile_23_clock; 
  wire  uRegFile_23_reset; 
  wire [31:0] uRegFile_23_io_q; 
  wire [31:0] uRegFile_23_io_d; 
  wire  uRegFile_23_io_clear; 
  wire  uRegFile_24_clock; 
  wire  uRegFile_24_reset; 
  wire [31:0] uRegFile_24_io_q; 
  wire [31:0] uRegFile_24_io_d; 
  wire  uRegFile_24_io_clear; 
  wire  uRegFile_25_clock; 
  wire  uRegFile_25_reset; 
  wire [31:0] uRegFile_25_io_q; 
  wire [31:0] uRegFile_25_io_d; 
  wire  uRegFile_25_io_clear; 
  wire  uRegFile_26_clock; 
  wire  uRegFile_26_reset; 
  wire [31:0] uRegFile_26_io_q; 
  wire [31:0] uRegFile_26_io_d; 
  wire  uRegFile_26_io_clear; 
  wire  uRegFile_27_clock; 
  wire  uRegFile_27_reset; 
  wire [31:0] uRegFile_27_io_q; 
  wire [31:0] uRegFile_27_io_d; 
  wire  uRegFile_27_io_clear; 
  wire  uRegFile_28_clock; 
  wire  uRegFile_28_reset; 
  wire [31:0] uRegFile_28_io_q; 
  wire [31:0] uRegFile_28_io_d; 
  wire  uRegFile_28_io_clear; 
  wire  uRegFile_29_clock; 
  wire  uRegFile_29_reset; 
  wire [31:0] uRegFile_29_io_q; 
  wire [31:0] uRegFile_29_io_d; 
  wire  uRegFile_29_io_clear; 
  wire  uRegFile_30_clock; 
  wire  uRegFile_30_reset; 
  wire [31:0] uRegFile_30_io_q; 
  wire [31:0] uRegFile_30_io_d; 
  wire  uRegFile_30_io_clear; 
  wire  uRegFile_31_clock; 
  wire  uRegFile_31_reset; 
  wire [31:0] uRegFile_31_io_q; 
  wire [31:0] uRegFile_31_io_d; 
  wire  uRegFile_31_io_clear; 
  wire  uRegState_0_clock; 
  wire  uRegState_0_reset; 
  wire  uRegState_0_io_q_busy; 
  wire [4:0] uRegState_0_io_q_reorder; 
  wire  uRegState_0_io_d_busy; 
  wire [4:0] uRegState_0_io_d_reorder; 
  wire  uRegState_0_io_clear; 
  wire  uRegState_1_clock; 
  wire  uRegState_1_reset; 
  wire  uRegState_1_io_q_busy; 
  wire [4:0] uRegState_1_io_q_reorder; 
  wire  uRegState_1_io_d_busy; 
  wire [4:0] uRegState_1_io_d_reorder; 
  wire  uRegState_1_io_clear; 
  wire  uRegState_2_clock; 
  wire  uRegState_2_reset; 
  wire  uRegState_2_io_q_busy; 
  wire [4:0] uRegState_2_io_q_reorder; 
  wire  uRegState_2_io_d_busy; 
  wire [4:0] uRegState_2_io_d_reorder; 
  wire  uRegState_2_io_clear; 
  wire  uRegState_3_clock; 
  wire  uRegState_3_reset; 
  wire  uRegState_3_io_q_busy; 
  wire [4:0] uRegState_3_io_q_reorder; 
  wire  uRegState_3_io_d_busy; 
  wire [4:0] uRegState_3_io_d_reorder; 
  wire  uRegState_3_io_clear; 
  wire  uRegState_4_clock; 
  wire  uRegState_4_reset; 
  wire  uRegState_4_io_q_busy; 
  wire [4:0] uRegState_4_io_q_reorder; 
  wire  uRegState_4_io_d_busy; 
  wire [4:0] uRegState_4_io_d_reorder; 
  wire  uRegState_4_io_clear; 
  wire  uRegState_5_clock; 
  wire  uRegState_5_reset; 
  wire  uRegState_5_io_q_busy; 
  wire [4:0] uRegState_5_io_q_reorder; 
  wire  uRegState_5_io_d_busy; 
  wire [4:0] uRegState_5_io_d_reorder; 
  wire  uRegState_5_io_clear; 
  wire  uRegState_6_clock; 
  wire  uRegState_6_reset; 
  wire  uRegState_6_io_q_busy; 
  wire [4:0] uRegState_6_io_q_reorder; 
  wire  uRegState_6_io_d_busy; 
  wire [4:0] uRegState_6_io_d_reorder; 
  wire  uRegState_6_io_clear; 
  wire  uRegState_7_clock; 
  wire  uRegState_7_reset; 
  wire  uRegState_7_io_q_busy; 
  wire [4:0] uRegState_7_io_q_reorder; 
  wire  uRegState_7_io_d_busy; 
  wire [4:0] uRegState_7_io_d_reorder; 
  wire  uRegState_7_io_clear; 
  wire  uRegState_8_clock; 
  wire  uRegState_8_reset; 
  wire  uRegState_8_io_q_busy; 
  wire [4:0] uRegState_8_io_q_reorder; 
  wire  uRegState_8_io_d_busy; 
  wire [4:0] uRegState_8_io_d_reorder; 
  wire  uRegState_8_io_clear; 
  wire  uRegState_9_clock; 
  wire  uRegState_9_reset; 
  wire  uRegState_9_io_q_busy; 
  wire [4:0] uRegState_9_io_q_reorder; 
  wire  uRegState_9_io_d_busy; 
  wire [4:0] uRegState_9_io_d_reorder; 
  wire  uRegState_9_io_clear; 
  wire  uRegState_10_clock; 
  wire  uRegState_10_reset; 
  wire  uRegState_10_io_q_busy; 
  wire [4:0] uRegState_10_io_q_reorder; 
  wire  uRegState_10_io_d_busy; 
  wire [4:0] uRegState_10_io_d_reorder; 
  wire  uRegState_10_io_clear; 
  wire  uRegState_11_clock; 
  wire  uRegState_11_reset; 
  wire  uRegState_11_io_q_busy; 
  wire [4:0] uRegState_11_io_q_reorder; 
  wire  uRegState_11_io_d_busy; 
  wire [4:0] uRegState_11_io_d_reorder; 
  wire  uRegState_11_io_clear; 
  wire  uRegState_12_clock; 
  wire  uRegState_12_reset; 
  wire  uRegState_12_io_q_busy; 
  wire [4:0] uRegState_12_io_q_reorder; 
  wire  uRegState_12_io_d_busy; 
  wire [4:0] uRegState_12_io_d_reorder; 
  wire  uRegState_12_io_clear; 
  wire  uRegState_13_clock; 
  wire  uRegState_13_reset; 
  wire  uRegState_13_io_q_busy; 
  wire [4:0] uRegState_13_io_q_reorder; 
  wire  uRegState_13_io_d_busy; 
  wire [4:0] uRegState_13_io_d_reorder; 
  wire  uRegState_13_io_clear; 
  wire  uRegState_14_clock; 
  wire  uRegState_14_reset; 
  wire  uRegState_14_io_q_busy; 
  wire [4:0] uRegState_14_io_q_reorder; 
  wire  uRegState_14_io_d_busy; 
  wire [4:0] uRegState_14_io_d_reorder; 
  wire  uRegState_14_io_clear; 
  wire  uRegState_15_clock; 
  wire  uRegState_15_reset; 
  wire  uRegState_15_io_q_busy; 
  wire [4:0] uRegState_15_io_q_reorder; 
  wire  uRegState_15_io_d_busy; 
  wire [4:0] uRegState_15_io_d_reorder; 
  wire  uRegState_15_io_clear; 
  wire  uRegState_16_clock; 
  wire  uRegState_16_reset; 
  wire  uRegState_16_io_q_busy; 
  wire [4:0] uRegState_16_io_q_reorder; 
  wire  uRegState_16_io_d_busy; 
  wire [4:0] uRegState_16_io_d_reorder; 
  wire  uRegState_16_io_clear; 
  wire  uRegState_17_clock; 
  wire  uRegState_17_reset; 
  wire  uRegState_17_io_q_busy; 
  wire [4:0] uRegState_17_io_q_reorder; 
  wire  uRegState_17_io_d_busy; 
  wire [4:0] uRegState_17_io_d_reorder; 
  wire  uRegState_17_io_clear; 
  wire  uRegState_18_clock; 
  wire  uRegState_18_reset; 
  wire  uRegState_18_io_q_busy; 
  wire [4:0] uRegState_18_io_q_reorder; 
  wire  uRegState_18_io_d_busy; 
  wire [4:0] uRegState_18_io_d_reorder; 
  wire  uRegState_18_io_clear; 
  wire  uRegState_19_clock; 
  wire  uRegState_19_reset; 
  wire  uRegState_19_io_q_busy; 
  wire [4:0] uRegState_19_io_q_reorder; 
  wire  uRegState_19_io_d_busy; 
  wire [4:0] uRegState_19_io_d_reorder; 
  wire  uRegState_19_io_clear; 
  wire  uRegState_20_clock; 
  wire  uRegState_20_reset; 
  wire  uRegState_20_io_q_busy; 
  wire [4:0] uRegState_20_io_q_reorder; 
  wire  uRegState_20_io_d_busy; 
  wire [4:0] uRegState_20_io_d_reorder; 
  wire  uRegState_20_io_clear; 
  wire  uRegState_21_clock; 
  wire  uRegState_21_reset; 
  wire  uRegState_21_io_q_busy; 
  wire [4:0] uRegState_21_io_q_reorder; 
  wire  uRegState_21_io_d_busy; 
  wire [4:0] uRegState_21_io_d_reorder; 
  wire  uRegState_21_io_clear; 
  wire  uRegState_22_clock; 
  wire  uRegState_22_reset; 
  wire  uRegState_22_io_q_busy; 
  wire [4:0] uRegState_22_io_q_reorder; 
  wire  uRegState_22_io_d_busy; 
  wire [4:0] uRegState_22_io_d_reorder; 
  wire  uRegState_22_io_clear; 
  wire  uRegState_23_clock; 
  wire  uRegState_23_reset; 
  wire  uRegState_23_io_q_busy; 
  wire [4:0] uRegState_23_io_q_reorder; 
  wire  uRegState_23_io_d_busy; 
  wire [4:0] uRegState_23_io_d_reorder; 
  wire  uRegState_23_io_clear; 
  wire  uRegState_24_clock; 
  wire  uRegState_24_reset; 
  wire  uRegState_24_io_q_busy; 
  wire [4:0] uRegState_24_io_q_reorder; 
  wire  uRegState_24_io_d_busy; 
  wire [4:0] uRegState_24_io_d_reorder; 
  wire  uRegState_24_io_clear; 
  wire  uRegState_25_clock; 
  wire  uRegState_25_reset; 
  wire  uRegState_25_io_q_busy; 
  wire [4:0] uRegState_25_io_q_reorder; 
  wire  uRegState_25_io_d_busy; 
  wire [4:0] uRegState_25_io_d_reorder; 
  wire  uRegState_25_io_clear; 
  wire  uRegState_26_clock; 
  wire  uRegState_26_reset; 
  wire  uRegState_26_io_q_busy; 
  wire [4:0] uRegState_26_io_q_reorder; 
  wire  uRegState_26_io_d_busy; 
  wire [4:0] uRegState_26_io_d_reorder; 
  wire  uRegState_26_io_clear; 
  wire  uRegState_27_clock; 
  wire  uRegState_27_reset; 
  wire  uRegState_27_io_q_busy; 
  wire [4:0] uRegState_27_io_q_reorder; 
  wire  uRegState_27_io_d_busy; 
  wire [4:0] uRegState_27_io_d_reorder; 
  wire  uRegState_27_io_clear; 
  wire  uRegState_28_clock; 
  wire  uRegState_28_reset; 
  wire  uRegState_28_io_q_busy; 
  wire [4:0] uRegState_28_io_q_reorder; 
  wire  uRegState_28_io_d_busy; 
  wire [4:0] uRegState_28_io_d_reorder; 
  wire  uRegState_28_io_clear; 
  wire  uRegState_29_clock; 
  wire  uRegState_29_reset; 
  wire  uRegState_29_io_q_busy; 
  wire [4:0] uRegState_29_io_q_reorder; 
  wire  uRegState_29_io_d_busy; 
  wire [4:0] uRegState_29_io_d_reorder; 
  wire  uRegState_29_io_clear; 
  wire  uRegState_30_clock; 
  wire  uRegState_30_reset; 
  wire  uRegState_30_io_q_busy; 
  wire [4:0] uRegState_30_io_q_reorder; 
  wire  uRegState_30_io_d_busy; 
  wire [4:0] uRegState_30_io_d_reorder; 
  wire  uRegState_30_io_clear; 
  wire  uRegState_31_clock; 
  wire  uRegState_31_reset; 
  wire  uRegState_31_io_q_busy; 
  wire [4:0] uRegState_31_io_q_reorder; 
  wire  uRegState_31_io_d_busy; 
  wire [4:0] uRegState_31_io_d_reorder; 
  wire  uRegState_31_io_clear; 
  wire  integer_inst_r_clock; 
  wire  integer_inst_r_reset; 
  wire  integer_inst_r_io_q; 
  wire  integer_inst_r_io_d; 
  wire  integer_inst_r_io_clear; 
  wire  branch_inst_r_clock; 
  wire  branch_inst_r_reset; 
  wire  branch_inst_r_io_q; 
  wire  branch_inst_r_io_d; 
  wire  branch_inst_r_io_clear; 
  wire  store_inst_r_clock; 
  wire  store_inst_r_reset; 
  wire  store_inst_r_io_q; 
  wire  store_inst_r_io_d; 
  wire  store_inst_r_io_clear; 
  wire  load_inst_r_clock; 
  wire  load_inst_r_reset; 
  wire  load_inst_r_io_q; 
  wire  load_inst_r_io_d; 
  wire  load_inst_r_io_clear; 
  wire  muldiv_inst_r_clock; 
  wire  muldiv_inst_r_reset; 
  wire  muldiv_inst_r_io_q; 
  wire  muldiv_inst_r_io_d; 
  wire  muldiv_inst_r_io_clear; 
  wire  mBranchProc_st_clock; 
  wire  mBranchProc_st_reset; 
  wire [1:0] mBranchProc_st_io_q; 
  wire [1:0] mBranchProc_st_io_d; 
  wire  mBranchProc_st_io_clear; 
  wire  re_jump_addr_r_clock; 
  wire  re_jump_addr_r_reset; 
  wire [31:0] re_jump_addr_r_io_q; 
  wire [31:0] re_jump_addr_r_io_d; 
  wire  re_jump_addr_r_io_clear; 
  wire  uIntBusGetData_st_clock; 
  wire  uIntBusGetData_st_reset; 
  wire  uIntBusGetData_st_io_q; 
  wire  uIntBusGetData_st_io_d; 
  wire  uIntBusGetData_st_io_clear; 
  wire  uMulDivBusGetData_st_clock; 
  wire  uMulDivBusGetData_st_reset; 
  wire  uMulDivBusGetData_st_io_q; 
  wire  uMulDivBusGetData_st_io_d; 
  wire  uMulDivBusGetData_st_io_clear; 
  wire  uLoadBusGetData_st_clock; 
  wire  uLoadBusGetData_st_reset; 
  wire  uLoadBusGetData_st_io_q; 
  wire  uLoadBusGetData_st_io_d; 
  wire  uLoadBusGetData_st_io_clear; 
  wire  uROB_io_queue_data_split_0_rob_ready = uROB__io_queue_data[0]; 
  wire [31:0] uROB_io_queue_data_split_0_rob_value = uROB__io_queue_data[32:1]; 
  wire  uROB_io_queue_data_split_1_rob_ready = uROB__io_queue_data[67]; 
  wire [31:0] uROB_io_queue_data_split_1_rob_value = uROB__io_queue_data[99:68]; 
  wire [31:0] uROB_io_queue_data_split_1_rob_dest = uROB__io_queue_data[131:100]; 
  wire [1:0] uROB_io_queue_data_split_1_rob_type = uROB__io_queue_data[133:132]; 
  wire  uROB_io_queue_data_split_2_rob_ready = uROB__io_queue_data[134]; 
  wire [31:0] uROB_io_queue_data_split_2_rob_value = uROB__io_queue_data[166:135]; 
  wire [31:0] uROB_io_queue_data_split_2_rob_dest = uROB__io_queue_data[198:167]; 
  wire [1:0] uROB_io_queue_data_split_2_rob_type = uROB__io_queue_data[200:199]; 
  wire  uROB_io_queue_data_split_3_rob_ready = uROB__io_queue_data[201]; 
  wire [31:0] uROB_io_queue_data_split_3_rob_value = uROB__io_queue_data[233:202]; 
  wire [31:0] uROB_io_queue_data_split_3_rob_dest = uROB__io_queue_data[265:234]; 
  wire [1:0] uROB_io_queue_data_split_3_rob_type = uROB__io_queue_data[267:266]; 
  wire  uROB_io_queue_data_split_4_rob_ready = uROB__io_queue_data[268]; 
  wire [31:0] uROB_io_queue_data_split_4_rob_value = uROB__io_queue_data[300:269]; 
  wire [31:0] uROB_io_queue_data_split_4_rob_dest = uROB__io_queue_data[332:301]; 
  wire [1:0] uROB_io_queue_data_split_4_rob_type = uROB__io_queue_data[334:333]; 
  wire  uROB_io_queue_data_split_5_rob_ready = uROB__io_queue_data[335]; 
  wire [31:0] uROB_io_queue_data_split_5_rob_value = uROB__io_queue_data[367:336]; 
  wire [31:0] uROB_io_queue_data_split_5_rob_dest = uROB__io_queue_data[399:368]; 
  wire [1:0] uROB_io_queue_data_split_5_rob_type = uROB__io_queue_data[401:400]; 
  wire  uROB_io_queue_data_split_6_rob_ready = uROB__io_queue_data[402]; 
  wire [31:0] uROB_io_queue_data_split_6_rob_value = uROB__io_queue_data[434:403]; 
  wire [31:0] uROB_io_queue_data_split_6_rob_dest = uROB__io_queue_data[466:435]; 
  wire [1:0] uROB_io_queue_data_split_6_rob_type = uROB__io_queue_data[468:467]; 
  wire  uROB_io_queue_data_split_7_rob_ready = uROB__io_queue_data[469]; 
  wire [31:0] uROB_io_queue_data_split_7_rob_value = uROB__io_queue_data[501:470]; 
  wire [31:0] uROB_io_queue_data_split_7_rob_dest = uROB__io_queue_data[533:502]; 
  wire [1:0] uROB_io_queue_data_split_7_rob_type = uROB__io_queue_data[535:534]; 
  wire  uROB_io_queue_data_split_8_rob_ready = uROB__io_queue_data[536]; 
  wire [31:0] uROB_io_queue_data_split_8_rob_value = uROB__io_queue_data[568:537]; 
  wire [31:0] uROB_io_queue_data_split_8_rob_dest = uROB__io_queue_data[600:569]; 
  wire [1:0] uROB_io_queue_data_split_8_rob_type = uROB__io_queue_data[602:601]; 
  wire  uROB_io_queue_data_split_9_rob_ready = uROB__io_queue_data[603]; 
  wire [31:0] uROB_io_queue_data_split_9_rob_value = uROB__io_queue_data[635:604]; 
  wire [31:0] uROB_io_queue_data_split_9_rob_dest = uROB__io_queue_data[667:636]; 
  wire [1:0] uROB_io_queue_data_split_9_rob_type = uROB__io_queue_data[669:668]; 
  wire  uROB_io_queue_data_split_10_rob_ready = uROB__io_queue_data[670]; 
  wire [31:0] uROB_io_queue_data_split_10_rob_value = uROB__io_queue_data[702:671]; 
  wire [31:0] uROB_io_queue_data_split_10_rob_dest = uROB__io_queue_data[734:703]; 
  wire [1:0] uROB_io_queue_data_split_10_rob_type = uROB__io_queue_data[736:735]; 
  wire  uROB_io_queue_data_split_11_rob_ready = uROB__io_queue_data[737]; 
  wire [31:0] uROB_io_queue_data_split_11_rob_value = uROB__io_queue_data[769:738]; 
  wire [31:0] uROB_io_queue_data_split_11_rob_dest = uROB__io_queue_data[801:770]; 
  wire [1:0] uROB_io_queue_data_split_11_rob_type = uROB__io_queue_data[803:802]; 
  wire  uROB_io_queue_data_split_12_rob_ready = uROB__io_queue_data[804]; 
  wire [31:0] uROB_io_queue_data_split_12_rob_value = uROB__io_queue_data[836:805]; 
  wire [31:0] uROB_io_queue_data_split_12_rob_dest = uROB__io_queue_data[868:837]; 
  wire [1:0] uROB_io_queue_data_split_12_rob_type = uROB__io_queue_data[870:869]; 
  wire  uROB_io_queue_data_split_13_rob_ready = uROB__io_queue_data[871]; 
  wire [31:0] uROB_io_queue_data_split_13_rob_value = uROB__io_queue_data[903:872]; 
  wire [31:0] uROB_io_queue_data_split_13_rob_dest = uROB__io_queue_data[935:904]; 
  wire [1:0] uROB_io_queue_data_split_13_rob_type = uROB__io_queue_data[937:936]; 
  wire  uROB_io_queue_data_split_14_rob_ready = uROB__io_queue_data[938]; 
  wire [31:0] uROB_io_queue_data_split_14_rob_value = uROB__io_queue_data[970:939]; 
  wire [31:0] uROB_io_queue_data_split_14_rob_dest = uROB__io_queue_data[1002:971]; 
  wire [1:0] uROB_io_queue_data_split_14_rob_type = uROB__io_queue_data[1004:1003]; 
  wire  uROB_io_queue_data_split_15_rob_ready = uROB__io_queue_data[1005]; 
  wire [31:0] uROB_io_queue_data_split_15_rob_value = uROB__io_queue_data[1037:1006]; 
  wire [31:0] uROB_io_queue_data_split_15_rob_dest = uROB__io_queue_data[1069:1038]; 
  wire [1:0] uROB_io_queue_data_split_15_rob_type = uROB__io_queue_data[1071:1070]; 
  wire  uROB_io_queue_data_split_16_rob_ready = uROB__io_queue_data[1072]; 
  wire [31:0] uROB_io_queue_data_split_16_rob_value = uROB__io_queue_data[1104:1073]; 
  wire [31:0] uROB_io_queue_data_split_16_rob_dest = uROB__io_queue_data[1136:1105]; 
  wire [1:0] uROB_io_queue_data_split_16_rob_type = uROB__io_queue_data[1138:1137]; 
  wire [19:0] uLoadStoreRS_io_deq_data_op = uLoadStoreRS__io_deq_data[131:112]; 
  wire  uLoadstoreRS_deq_data_op_store = uLoadStoreRS_io_deq_data_op[19]; 
  wire [4:0] uLoadStoreRS_io_deq_data_qj = uLoadStoreRS__io_deq_data[106:102]; 
  wire  _uLoadStoreRS_out_valid_T_1 = uLoadStoreRS_io_deq_data_qj == 5'h0; 
  wire  _uLoadStoreRS_out_valid_T_2 = ~uLoadStoreRS__io_empty & _uLoadStoreRS_out_valid_T_1; 
  wire [4:0] uLoadStoreRS_io_deq_data_qk = uLoadStoreRS__io_deq_data[101:97]; 
  wire  _uLoadStoreRS_out_valid_T_3 = uLoadStoreRS_io_deq_data_qk == 5'h0; 
  wire  uLoadStoreRS_out_valid = _uLoadStoreRS_out_valid_T_2 & _uLoadStoreRS_out_valid_T_3; 
  wire  set_ROB_store_ready = uLoadstoreRS_deq_data_op_store & uLoadStoreRS_out_valid; 
  wire [4:0] uLoadStoreRS_io_deq_data_dest = uLoadStoreRS__io_deq_data[111:107]; 
  wire  _T_428 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h1; 
  wire [31:0] uLoadStoreRS_io_deq_data_vk = uLoadStoreRS__io_deq_data[32:1]; 
  wire [31:0] _GEN_2601 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h1 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_1_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_1_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h1 ?
    uCDB_io_cdb_result : _GEN_2601; 
  wire  _GEN_2602 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h1 | uROB_io_queue_data_split_1_rob_ready; 
  wire  uROB_io_update_entry_data_split_1_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h1 | _GEN_2602; 
  wire [31:0] uLoadStoreRS_io_deq_data_vj = uLoadStoreRS__io_deq_data[64:33]; 
  wire [31:0] uLoadStoreRS_io_deq_data_a = uLoadStoreRS__io_deq_data[96:65]; 
  wire [31:0] issue_mem_addr = uLoadStoreRS_io_deq_data_vj + uLoadStoreRS_io_deq_data_a; 
  wire [31:0] _GEN_2600 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h1 ? issue_mem_addr :
    uROB_io_queue_data_split_1_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_1_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h1 ?
    uROB_io_queue_data_split_1_rob_dest : _GEN_2600; 
  wire [133:0] uROB_io_update_entry_data_lo_lo_lo = {uROB_io_queue_data_split_1_rob_type,
    uROB_io_update_entry_data_split_1_rob_dest,uROB_io_update_entry_data_split_1_rob_value,
    uROB_io_update_entry_data_split_1_rob_ready,67'h0}; 
  wire  _T_434 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h2; 
  wire [31:0] _GEN_2611 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h2 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_2_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_2_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h2 ?
    uCDB_io_cdb_result : _GEN_2611; 
  wire  _GEN_2612 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h2 | uROB_io_queue_data_split_2_rob_ready; 
  wire  uROB_io_update_entry_data_split_2_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h2 | _GEN_2612; 
  wire [31:0] _GEN_2610 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h2 ? issue_mem_addr :
    uROB_io_queue_data_split_2_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_2_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h2 ?
    uROB_io_queue_data_split_2_rob_dest : _GEN_2610; 
  wire  _T_440 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h3; 
  wire [31:0] _GEN_2621 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h3 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_3_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_3_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h3 ?
    uCDB_io_cdb_result : _GEN_2621; 
  wire  _GEN_2622 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h3 | uROB_io_queue_data_split_3_rob_ready; 
  wire  uROB_io_update_entry_data_split_3_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h3 | _GEN_2622; 
  wire  _T_446 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h4; 
  wire  _GEN_2632 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h4 | uROB_io_queue_data_split_4_rob_ready; 
  wire  uROB_io_update_entry_data_split_4_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h4 | _GEN_2632; 
  wire [31:0] _GEN_2620 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h3 ? issue_mem_addr :
    uROB_io_queue_data_split_3_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_3_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h3 ?
    uROB_io_queue_data_split_3_rob_dest : _GEN_2620; 
  wire [268:0] uROB_io_update_entry_data_lo_lo = {uROB_io_update_entry_data_split_4_rob_ready,
    uROB_io_queue_data_split_3_rob_type,uROB_io_update_entry_data_split_3_rob_dest,
    uROB_io_update_entry_data_split_3_rob_value,uROB_io_update_entry_data_split_3_rob_ready,
    uROB_io_queue_data_split_2_rob_type,uROB_io_update_entry_data_split_2_rob_dest,
    uROB_io_update_entry_data_split_2_rob_value,uROB_io_update_entry_data_split_2_rob_ready,
    uROB_io_update_entry_data_lo_lo_lo}; 
  wire [31:0] _GEN_2630 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h4 ? issue_mem_addr :
    uROB_io_queue_data_split_4_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_4_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h4 ?
    uROB_io_queue_data_split_4_rob_dest : _GEN_2630; 
  wire [31:0] _GEN_2631 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h4 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_4_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_4_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h4 ?
    uCDB_io_cdb_result : _GEN_2631; 
  wire  _T_452 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h5; 
  wire  _GEN_2642 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h5 | uROB_io_queue_data_split_5_rob_ready; 
  wire  uROB_io_update_entry_data_split_5_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h5 | _GEN_2642; 
  wire [31:0] _GEN_2640 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h5 ? issue_mem_addr :
    uROB_io_queue_data_split_5_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_5_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h5 ?
    uROB_io_queue_data_split_5_rob_dest : _GEN_2640; 
  wire [31:0] _GEN_2641 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h5 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_5_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_5_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h5 ?
    uCDB_io_cdb_result : _GEN_2641; 
  wire  _T_458 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h6; 
  wire  _GEN_2652 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h6 | uROB_io_queue_data_split_6_rob_ready; 
  wire  uROB_io_update_entry_data_split_6_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h6 | _GEN_2652; 
  wire [133:0] uROB_io_update_entry_data_lo_hi_lo = {uROB_io_update_entry_data_split_6_rob_ready,
    uROB_io_queue_data_split_5_rob_type,uROB_io_update_entry_data_split_5_rob_dest,
    uROB_io_update_entry_data_split_5_rob_value,uROB_io_update_entry_data_split_5_rob_ready,
    uROB_io_queue_data_split_4_rob_type,uROB_io_update_entry_data_split_4_rob_dest,
    uROB_io_update_entry_data_split_4_rob_value}; 
  wire [31:0] _GEN_2650 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h6 ? issue_mem_addr :
    uROB_io_queue_data_split_6_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_6_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h6 ?
    uROB_io_queue_data_split_6_rob_dest : _GEN_2650; 
  wire [31:0] _GEN_2651 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h6 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_6_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_6_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h6 ?
    uCDB_io_cdb_result : _GEN_2651; 
  wire  _T_464 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h7; 
  wire  _GEN_2662 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h7 | uROB_io_queue_data_split_7_rob_ready; 
  wire  uROB_io_update_entry_data_split_7_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h7 | _GEN_2662; 
  wire [31:0] _GEN_2660 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h7 ? issue_mem_addr :
    uROB_io_queue_data_split_7_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_7_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h7 ?
    uROB_io_queue_data_split_7_rob_dest : _GEN_2660; 
  wire [31:0] _GEN_2661 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h7 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_7_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_7_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h7 ?
    uCDB_io_cdb_result : _GEN_2661; 
  wire  _T_470 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h8; 
  wire [31:0] _GEN_2671 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h8 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_8_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_8_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h8 ?
    uCDB_io_cdb_result : _GEN_2671; 
  wire  _GEN_2672 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h8 | uROB_io_queue_data_split_8_rob_ready; 
  wire  uROB_io_update_entry_data_split_8_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h8 | _GEN_2672; 
  wire [299:0] uROB_io_update_entry_data_lo_hi = {uROB_io_update_entry_data_split_8_rob_value,
    uROB_io_update_entry_data_split_8_rob_ready,uROB_io_queue_data_split_7_rob_type,
    uROB_io_update_entry_data_split_7_rob_dest,uROB_io_update_entry_data_split_7_rob_value,
    uROB_io_update_entry_data_split_7_rob_ready,uROB_io_queue_data_split_6_rob_type,
    uROB_io_update_entry_data_split_6_rob_dest,uROB_io_update_entry_data_split_6_rob_value,
    uROB_io_update_entry_data_lo_hi_lo}; 
  wire [568:0] uROB_io_update_entry_data_lo = {uROB_io_update_entry_data_lo_hi,uROB_io_update_entry_data_lo_lo}; 
  wire [31:0] _GEN_2670 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h8 ? issue_mem_addr :
    uROB_io_queue_data_split_8_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_8_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h8 ?
    uROB_io_queue_data_split_8_rob_dest : _GEN_2670; 
  wire  _T_476 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h9; 
  wire [31:0] _GEN_2681 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h9 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_9_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_9_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h9 ?
    uCDB_io_cdb_result : _GEN_2681; 
  wire  _GEN_2682 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h9 | uROB_io_queue_data_split_9_rob_ready; 
  wire  uROB_io_update_entry_data_split_9_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h9 | _GEN_2682; 
  wire [31:0] _GEN_2680 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h9 ? issue_mem_addr :
    uROB_io_queue_data_split_9_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_9_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h9 ?
    uROB_io_queue_data_split_9_rob_dest : _GEN_2680; 
  wire  _T_482 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'ha; 
  wire [31:0] _GEN_2691 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'ha ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_10_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_10_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'ha ?
    uCDB_io_cdb_result : _GEN_2691; 
  wire  _GEN_2692 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'ha | uROB_io_queue_data_split_10_rob_ready; 
  wire  uROB_io_update_entry_data_split_10_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'ha | _GEN_2692; 
  wire [133:0] uROB_io_update_entry_data_hi_lo_lo = {uROB_io_update_entry_data_split_10_rob_value,
    uROB_io_update_entry_data_split_10_rob_ready,uROB_io_queue_data_split_9_rob_type,
    uROB_io_update_entry_data_split_9_rob_dest,uROB_io_update_entry_data_split_9_rob_value,
    uROB_io_update_entry_data_split_9_rob_ready,uROB_io_queue_data_split_8_rob_type,
    uROB_io_update_entry_data_split_8_rob_dest}; 
  wire [31:0] _GEN_2690 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'ha ? issue_mem_addr :
    uROB_io_queue_data_split_10_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_10_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'ha ?
    uROB_io_queue_data_split_10_rob_dest : _GEN_2690; 
  wire  _T_488 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hb; 
  wire [31:0] _GEN_2701 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hb ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_11_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_11_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hb ?
    uCDB_io_cdb_result : _GEN_2701; 
  wire  _GEN_2702 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hb | uROB_io_queue_data_split_11_rob_ready; 
  wire  uROB_io_update_entry_data_split_11_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hb | _GEN_2702; 
  wire [31:0] _GEN_2700 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hb ? issue_mem_addr :
    uROB_io_queue_data_split_11_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_11_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hb ?
    uROB_io_queue_data_split_11_rob_dest : _GEN_2700; 
  wire  _T_494 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hc; 
  wire [31:0] _GEN_2710 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hc ? issue_mem_addr :
    uROB_io_queue_data_split_12_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_12_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hc ?
    uROB_io_queue_data_split_12_rob_dest : _GEN_2710; 
  wire [31:0] _GEN_2711 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hc ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_12_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_12_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hc ?
    uCDB_io_cdb_result : _GEN_2711; 
  wire  _GEN_2712 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hc | uROB_io_queue_data_split_12_rob_ready; 
  wire  uROB_io_update_entry_data_split_12_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hc | _GEN_2712; 
  wire [299:0] uROB_io_update_entry_data_hi_lo = {uROB_io_update_entry_data_split_12_rob_dest,
    uROB_io_update_entry_data_split_12_rob_value,uROB_io_update_entry_data_split_12_rob_ready,
    uROB_io_queue_data_split_11_rob_type,uROB_io_update_entry_data_split_11_rob_dest,
    uROB_io_update_entry_data_split_11_rob_value,uROB_io_update_entry_data_split_11_rob_ready,
    uROB_io_queue_data_split_10_rob_type,uROB_io_update_entry_data_split_10_rob_dest,uROB_io_update_entry_data_hi_lo_lo}
    ; 
  wire  _T_500 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hd; 
  wire  _GEN_2722 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hd | uROB_io_queue_data_split_13_rob_ready; 
  wire  uROB_io_update_entry_data_split_13_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hd | _GEN_2722; 
  wire [31:0] _GEN_2720 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hd ? issue_mem_addr :
    uROB_io_queue_data_split_13_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_13_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hd ?
    uROB_io_queue_data_split_13_rob_dest : _GEN_2720; 
  wire [31:0] _GEN_2721 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hd ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_13_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_13_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hd ?
    uCDB_io_cdb_result : _GEN_2721; 
  wire  _T_506 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'he; 
  wire  _GEN_2732 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'he | uROB_io_queue_data_split_14_rob_ready; 
  wire  uROB_io_update_entry_data_split_14_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'he | _GEN_2732; 
  wire [31:0] _GEN_2730 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'he ? issue_mem_addr :
    uROB_io_queue_data_split_14_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_14_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'he ?
    uROB_io_queue_data_split_14_rob_dest : _GEN_2730; 
  wire [31:0] _GEN_2731 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'he ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_14_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_14_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'he ?
    uCDB_io_cdb_result : _GEN_2731; 
  wire [133:0] uROB_io_update_entry_data_hi_hi_lo = {uROB_io_update_entry_data_split_14_rob_dest,
    uROB_io_update_entry_data_split_14_rob_value,uROB_io_update_entry_data_split_14_rob_ready,
    uROB_io_queue_data_split_13_rob_type,uROB_io_update_entry_data_split_13_rob_dest,
    uROB_io_update_entry_data_split_13_rob_value,uROB_io_update_entry_data_split_13_rob_ready,
    uROB_io_queue_data_split_12_rob_type}; 
  wire  _T_512 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hf; 
  wire  _GEN_2742 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hf | uROB_io_queue_data_split_15_rob_ready; 
  wire  uROB_io_update_entry_data_split_15_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hf | _GEN_2742; 
  wire [31:0] _GEN_2740 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hf ? issue_mem_addr :
    uROB_io_queue_data_split_15_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_15_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hf ?
    uROB_io_queue_data_split_15_rob_dest : _GEN_2740; 
  wire [31:0] _GEN_2741 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'hf ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_15_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_15_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hf ?
    uCDB_io_cdb_result : _GEN_2741; 
  wire  _T_518 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h10; 
  wire  _GEN_2752 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h10 | uROB_io_queue_data_split_16_rob_ready
    ; 
  wire  uROB_io_update_entry_data_split_16_rob_ready = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h10 | _GEN_2752; 
  wire [31:0] _GEN_2750 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h10 ? issue_mem_addr :
    uROB_io_queue_data_split_16_rob_dest; 
  wire [31:0] uROB_io_update_entry_data_split_16_rob_dest = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h10 ?
    uROB_io_queue_data_split_16_rob_dest : _GEN_2750; 
  wire [31:0] _GEN_2751 = set_ROB_store_ready & uLoadStoreRS_io_deq_data_dest == 5'h10 ? uLoadStoreRS_io_deq_data_vk :
    uROB_io_queue_data_split_16_rob_value; 
  wire [31:0] uROB_io_update_entry_data_split_16_rob_value = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h10 ?
    uCDB_io_cdb_result : _GEN_2751; 
  wire [269:0] uROB_io_update_entry_data_hi_hi = {uROB_io_queue_data_split_16_rob_type,
    uROB_io_update_entry_data_split_16_rob_dest,uROB_io_update_entry_data_split_16_rob_value,
    uROB_io_update_entry_data_split_16_rob_ready,uROB_io_queue_data_split_15_rob_type,
    uROB_io_update_entry_data_split_15_rob_dest,uROB_io_update_entry_data_split_15_rob_value,
    uROB_io_update_entry_data_split_15_rob_ready,uROB_io_queue_data_split_14_rob_type,uROB_io_update_entry_data_hi_hi_lo
    }; 
  wire [569:0] uROB_io_update_entry_data_hi = {uROB_io_update_entry_data_hi_hi,uROB_io_update_entry_data_hi_lo}; 
  wire  uROB_io_update_entry_1 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h1 | _T_428; 
  wire  uROB_io_update_entry_3 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h3 | _T_440; 
  wire  uROB_io_update_entry_2 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h2 | _T_434; 
  wire  uROB_io_update_entry_5 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h5 | _T_452; 
  wire  uROB_io_update_entry_4 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h4 | _T_446; 
  wire  uROB_io_update_entry_7 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h7 | _T_464; 
  wire  uROB_io_update_entry_6 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h6 | _T_458; 
  wire [7:0] uROB_io_update_entry_lo = {uROB_io_update_entry_7,uROB_io_update_entry_6,uROB_io_update_entry_5,
    uROB_io_update_entry_4,uROB_io_update_entry_3,uROB_io_update_entry_2,uROB_io_update_entry_1,1'h0}; 
  wire  uROB_io_update_entry_9 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h9 | _T_476; 
  wire  uROB_io_update_entry_8 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h8 | _T_470; 
  wire  uROB_io_update_entry_11 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hb | _T_488; 
  wire  uROB_io_update_entry_10 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'ha | _T_482; 
  wire  uROB_io_update_entry_13 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hd | _T_500; 
  wire  uROB_io_update_entry_12 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hc | _T_494; 
  wire  uROB_io_update_entry_16 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'h10 | _T_518; 
  wire  uROB_io_update_entry_15 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'hf | _T_512; 
  wire  uROB_io_update_entry_14 = uCDB_io_cdb_valid & uCDB_io_cdb_dest == 5'he | _T_506; 
  wire [8:0] uROB_io_update_entry_hi = {uROB_io_update_entry_16,uROB_io_update_entry_15,uROB_io_update_entry_14,
    uROB_io_update_entry_13,uROB_io_update_entry_12,uROB_io_update_entry_11,uROB_io_update_entry_10,
    uROB_io_update_entry_9,uROB_io_update_entry_8}; 
  wire  _T_351 = ~uROB__io_full; 
  wire  _T_352 = ~uIntergerRS__io_full & ~uROB__io_full; 
  wire  _T_384 = ~uLoadStoreRS__io_full & _T_351; 
  wire  _T_406 = muldiv_inst_r_io_d; 
  wire  _T_409 = ~uMulDivRS__io_full & _T_351; 
  wire [1:0] _GEN_492 = ~uIntergerRS__io_full & ~uROB__io_full ? 2'h1 : 2'h0; 
  wire [1:0] _GEN_906 = _T_352 ? 2'h2 : 2'h0; 
  wire [1:0] _GEN_1256 = ~uLoadStoreRS__io_full & _T_351 ? 2'h3 : 2'h0; 
  wire [1:0] _GEN_1533 = _T_384 ? 2'h1 : 2'h0; 
  wire [1:0] _GEN_2012 = ~uMulDivRS__io_full & _T_351 ? 2'h1 : 2'h0; 
  wire [1:0] _GEN_2086 = muldiv_inst_r_io_d ? _GEN_2012 : 2'h0; 
  wire [1:0] _GEN_2160 = load_inst_r_io_d ? _GEN_1533 : _GEN_2086; 
  wire [1:0] _GEN_2243 = store_inst_r_io_d ? _GEN_1256 : _GEN_2160; 
  wire [1:0] _GEN_2326 = branch_inst_r_io_d ? _GEN_906 : _GEN_2243; 
  wire [1:0] _GEN_2416 = integer_inst_r_io_d ? _GEN_492 : _GEN_2326; 
  wire [1:0] uROB_io_enq_data_rob_type = decoder_if_inst_valid ? _GEN_2416 : 2'h0; 
  wire [31:0] _GEN_493 = ~uIntergerRS__io_full & ~uROB__io_full ? {{27'd0}, decoder_if_rd_idx} : 32'h0; 
  wire [31:0] _uROB_io_enq_data_rob_dest_T_1 = decoder_if_pc_out + 32'h4; 
  wire [31:0] _GEN_907 = _T_352 ? _uROB_io_enq_data_rob_dest_T_1 : 32'h0; 
  wire [31:0] _GEN_1534 = _T_384 ? {{27'd0}, decoder_if_rd_idx} : 32'h0; 
  wire [31:0] _GEN_2013 = ~uMulDivRS__io_full & _T_351 ? {{27'd0}, decoder_if_rd_idx} : 32'h0; 
  wire [31:0] _GEN_2087 = muldiv_inst_r_io_d ? _GEN_2013 : 32'h0; 
  wire [31:0] _GEN_2161 = load_inst_r_io_d ? _GEN_1534 : _GEN_2087; 
  wire [31:0] _GEN_2244 = store_inst_r_io_d ? 32'h0 : _GEN_2161; 
  wire [31:0] _GEN_2327 = branch_inst_r_io_d ? _GEN_907 : _GEN_2244; 
  wire [31:0] _GEN_2417 = integer_inst_r_io_d ? _GEN_493 : _GEN_2327; 
  wire [31:0] uROB_io_enq_data_rob_dest = decoder_if_inst_valid ? _GEN_2417 : 32'h0; 
  wire [33:0] uROB_io_enq_data_hi = {uROB_io_enq_data_rob_type,uROB_io_enq_data_rob_dest}; 
  wire  uROB_io_deq_data_rob_ready = uROB__io_deq_data[0]; 
  wire [31:0] uROB_io_deq_data_rob_value = uROB__io_deq_data[32:1]; 
  wire [31:0] uROB_io_deq_data_rob_dest = uROB__io_deq_data[64:33]; 
  wire [1:0] uROB_io_deq_data_rob_type = uROB__io_deq_data[66:65]; 
  wire  uIntergerRS_io_queue_data_split_0_busy = uIntergerRS__io_queue_data[0]; 
  wire [31:0] uIntergerRS_io_queue_data_split_0_vk = uIntergerRS__io_queue_data[32:1]; 
  wire [31:0] uIntergerRS_io_queue_data_split_0_vj = uIntergerRS__io_queue_data[64:33]; 
  wire [31:0] uIntergerRS_io_queue_data_split_0_a = uIntergerRS__io_queue_data[96:65]; 
  wire [4:0] uIntergerRS_io_queue_data_split_0_qk = uIntergerRS__io_queue_data[101:97]; 
  wire [4:0] uIntergerRS_io_queue_data_split_0_qj = uIntergerRS__io_queue_data[106:102]; 
  wire [4:0] uIntergerRS_io_queue_data_split_0_dest = uIntergerRS__io_queue_data[111:107]; 
  wire [19:0] uIntergerRS_io_queue_data_split_0_op = uIntergerRS__io_queue_data[131:112]; 
  wire  uIntergerRS_io_queue_data_split_1_busy = uIntergerRS__io_queue_data[132]; 
  wire [31:0] uIntergerRS_io_queue_data_split_1_vk = uIntergerRS__io_queue_data[164:133]; 
  wire [31:0] uIntergerRS_io_queue_data_split_1_vj = uIntergerRS__io_queue_data[196:165]; 
  wire [31:0] uIntergerRS_io_queue_data_split_1_a = uIntergerRS__io_queue_data[228:197]; 
  wire [4:0] uIntergerRS_io_queue_data_split_1_qk = uIntergerRS__io_queue_data[233:229]; 
  wire [4:0] uIntergerRS_io_queue_data_split_1_qj = uIntergerRS__io_queue_data[238:234]; 
  wire [4:0] uIntergerRS_io_queue_data_split_1_dest = uIntergerRS__io_queue_data[243:239]; 
  wire [19:0] uIntergerRS_io_queue_data_split_1_op = uIntergerRS__io_queue_data[263:244]; 
  wire  uIntergerRS_io_queue_data_split_2_busy = uIntergerRS__io_queue_data[264]; 
  wire [31:0] uIntergerRS_io_queue_data_split_2_vk = uIntergerRS__io_queue_data[296:265]; 
  wire [31:0] uIntergerRS_io_queue_data_split_2_vj = uIntergerRS__io_queue_data[328:297]; 
  wire [31:0] uIntergerRS_io_queue_data_split_2_a = uIntergerRS__io_queue_data[360:329]; 
  wire [4:0] uIntergerRS_io_queue_data_split_2_qk = uIntergerRS__io_queue_data[365:361]; 
  wire [4:0] uIntergerRS_io_queue_data_split_2_qj = uIntergerRS__io_queue_data[370:366]; 
  wire [4:0] uIntergerRS_io_queue_data_split_2_dest = uIntergerRS__io_queue_data[375:371]; 
  wire [19:0] uIntergerRS_io_queue_data_split_2_op = uIntergerRS__io_queue_data[395:376]; 
  wire  uIntergerRS_io_queue_data_split_3_busy = uIntergerRS__io_queue_data[396]; 
  wire [31:0] uIntergerRS_io_queue_data_split_3_vk = uIntergerRS__io_queue_data[428:397]; 
  wire [31:0] uIntergerRS_io_queue_data_split_3_vj = uIntergerRS__io_queue_data[460:429]; 
  wire [31:0] uIntergerRS_io_queue_data_split_3_a = uIntergerRS__io_queue_data[492:461]; 
  wire [4:0] uIntergerRS_io_queue_data_split_3_qk = uIntergerRS__io_queue_data[497:493]; 
  wire [4:0] uIntergerRS_io_queue_data_split_3_qj = uIntergerRS__io_queue_data[502:498]; 
  wire [4:0] uIntergerRS_io_queue_data_split_3_dest = uIntergerRS__io_queue_data[507:503]; 
  wire [19:0] uIntergerRS_io_queue_data_split_3_op = uIntergerRS__io_queue_data[527:508]; 
  wire  uRegState_io_31_q_busy = uRegState_31_io_q_busy; 
  wire  uRegState_io_30_q_busy = uRegState_30_io_q_busy; 
  wire  uRegState_io_29_q_busy = uRegState_29_io_q_busy; 
  wire  uRegState_io_28_q_busy = uRegState_28_io_q_busy; 
  wire  uRegState_io_27_q_busy = uRegState_27_io_q_busy; 
  wire  uRegState_io_26_q_busy = uRegState_26_io_q_busy; 
  wire  uRegState_io_25_q_busy = uRegState_25_io_q_busy; 
  wire  uRegState_io_24_q_busy = uRegState_24_io_q_busy; 
  wire  uRegState_io_23_q_busy = uRegState_23_io_q_busy; 
  wire  uRegState_io_22_q_busy = uRegState_22_io_q_busy; 
  wire  uRegState_io_21_q_busy = uRegState_21_io_q_busy; 
  wire  uRegState_io_20_q_busy = uRegState_20_io_q_busy; 
  wire  uRegState_io_19_q_busy = uRegState_19_io_q_busy; 
  wire  uRegState_io_18_q_busy = uRegState_18_io_q_busy; 
  wire  uRegState_io_17_q_busy = uRegState_17_io_q_busy; 
  wire  uRegState_io_16_q_busy = uRegState_16_io_q_busy; 
  wire  uRegState_io_15_q_busy = uRegState_15_io_q_busy; 
  wire  uRegState_io_14_q_busy = uRegState_14_io_q_busy; 
  wire  uRegState_io_13_q_busy = uRegState_13_io_q_busy; 
  wire  uRegState_io_12_q_busy = uRegState_12_io_q_busy; 
  wire  uRegState_io_11_q_busy = uRegState_11_io_q_busy; 
  wire  uRegState_io_10_q_busy = uRegState_10_io_q_busy; 
  wire  uRegState_io_9_q_busy = uRegState_9_io_q_busy; 
  wire  uRegState_io_8_q_busy = uRegState_8_io_q_busy; 
  wire  uRegState_io_7_q_busy = uRegState_7_io_q_busy; 
  wire  uRegState_io_6_q_busy = uRegState_6_io_q_busy; 
  wire  uRegState_io_5_q_busy = uRegState_5_io_q_busy; 
  wire  uRegState_io_4_q_busy = uRegState_4_io_q_busy; 
  wire  uRegState_io_3_q_busy = uRegState_3_io_q_busy; 
  wire  uRegState_io_2_q_busy = uRegState_2_io_q_busy; 
  wire  uRegState_io_1_q_busy = uRegState_1_io_q_busy; 
  wire  uRegState_io_0_q_busy = uRegState_0_io_q_busy; 
  wire  _GEN_355 = 5'h1 == decoder_if_rt_idx ? uRegState_io_1_q_busy : uRegState_io_0_q_busy; 
  wire  _GEN_356 = 5'h2 == decoder_if_rt_idx ? uRegState_io_2_q_busy : _GEN_355; 
  wire  _GEN_357 = 5'h3 == decoder_if_rt_idx ? uRegState_io_3_q_busy : _GEN_356; 
  wire  _GEN_358 = 5'h4 == decoder_if_rt_idx ? uRegState_io_4_q_busy : _GEN_357; 
  wire  _GEN_359 = 5'h5 == decoder_if_rt_idx ? uRegState_io_5_q_busy : _GEN_358; 
  wire  _GEN_360 = 5'h6 == decoder_if_rt_idx ? uRegState_io_6_q_busy : _GEN_359; 
  wire  _GEN_361 = 5'h7 == decoder_if_rt_idx ? uRegState_io_7_q_busy : _GEN_360; 
  wire  _GEN_362 = 5'h8 == decoder_if_rt_idx ? uRegState_io_8_q_busy : _GEN_361; 
  wire  _GEN_363 = 5'h9 == decoder_if_rt_idx ? uRegState_io_9_q_busy : _GEN_362; 
  wire  _GEN_364 = 5'ha == decoder_if_rt_idx ? uRegState_io_10_q_busy : _GEN_363; 
  wire  _GEN_365 = 5'hb == decoder_if_rt_idx ? uRegState_io_11_q_busy : _GEN_364; 
  wire  _GEN_366 = 5'hc == decoder_if_rt_idx ? uRegState_io_12_q_busy : _GEN_365; 
  wire  _GEN_367 = 5'hd == decoder_if_rt_idx ? uRegState_io_13_q_busy : _GEN_366; 
  wire  _GEN_368 = 5'he == decoder_if_rt_idx ? uRegState_io_14_q_busy : _GEN_367; 
  wire  _GEN_369 = 5'hf == decoder_if_rt_idx ? uRegState_io_15_q_busy : _GEN_368; 
  wire  _GEN_370 = 5'h10 == decoder_if_rt_idx ? uRegState_io_16_q_busy : _GEN_369; 
  wire  _GEN_371 = 5'h11 == decoder_if_rt_idx ? uRegState_io_17_q_busy : _GEN_370; 
  wire  _GEN_372 = 5'h12 == decoder_if_rt_idx ? uRegState_io_18_q_busy : _GEN_371; 
  wire  _GEN_373 = 5'h13 == decoder_if_rt_idx ? uRegState_io_19_q_busy : _GEN_372; 
  wire  _GEN_374 = 5'h14 == decoder_if_rt_idx ? uRegState_io_20_q_busy : _GEN_373; 
  wire  _GEN_375 = 5'h15 == decoder_if_rt_idx ? uRegState_io_21_q_busy : _GEN_374; 
  wire  _GEN_376 = 5'h16 == decoder_if_rt_idx ? uRegState_io_22_q_busy : _GEN_375; 
  wire  _GEN_377 = 5'h17 == decoder_if_rt_idx ? uRegState_io_23_q_busy : _GEN_376; 
  wire  _GEN_378 = 5'h18 == decoder_if_rt_idx ? uRegState_io_24_q_busy : _GEN_377; 
  wire  _GEN_379 = 5'h19 == decoder_if_rt_idx ? uRegState_io_25_q_busy : _GEN_378; 
  wire  _GEN_380 = 5'h1a == decoder_if_rt_idx ? uRegState_io_26_q_busy : _GEN_379; 
  wire  _GEN_381 = 5'h1b == decoder_if_rt_idx ? uRegState_io_27_q_busy : _GEN_380; 
  wire  _GEN_382 = 5'h1c == decoder_if_rt_idx ? uRegState_io_28_q_busy : _GEN_381; 
  wire  _GEN_383 = 5'h1d == decoder_if_rt_idx ? uRegState_io_29_q_busy : _GEN_382; 
  wire  _GEN_384 = 5'h1e == decoder_if_rt_idx ? uRegState_io_30_q_busy : _GEN_383; 
  wire  _GEN_385 = 5'h1f == decoder_if_rt_idx ? uRegState_io_31_q_busy : _GEN_384; 
  wire [4:0] uRegState_io_31_q_reorder = uRegState_31_io_q_reorder; 
  wire [4:0] uRegState_io_30_q_reorder = uRegState_30_io_q_reorder; 
  wire [4:0] uRegState_io_29_q_reorder = uRegState_29_io_q_reorder; 
  wire [4:0] uRegState_io_28_q_reorder = uRegState_28_io_q_reorder; 
  wire [4:0] uRegState_io_27_q_reorder = uRegState_27_io_q_reorder; 
  wire [4:0] uRegState_io_26_q_reorder = uRegState_26_io_q_reorder; 
  wire [4:0] uRegState_io_25_q_reorder = uRegState_25_io_q_reorder; 
  wire [4:0] uRegState_io_24_q_reorder = uRegState_24_io_q_reorder; 
  wire [4:0] uRegState_io_23_q_reorder = uRegState_23_io_q_reorder; 
  wire [4:0] uRegState_io_22_q_reorder = uRegState_22_io_q_reorder; 
  wire [4:0] uRegState_io_21_q_reorder = uRegState_21_io_q_reorder; 
  wire [4:0] uRegState_io_20_q_reorder = uRegState_20_io_q_reorder; 
  wire [4:0] uRegState_io_19_q_reorder = uRegState_19_io_q_reorder; 
  wire [4:0] uRegState_io_18_q_reorder = uRegState_18_io_q_reorder; 
  wire [4:0] uRegState_io_17_q_reorder = uRegState_17_io_q_reorder; 
  wire [4:0] uRegState_io_16_q_reorder = uRegState_16_io_q_reorder; 
  wire [4:0] uRegState_io_15_q_reorder = uRegState_15_io_q_reorder; 
  wire [4:0] uRegState_io_14_q_reorder = uRegState_14_io_q_reorder; 
  wire [4:0] uRegState_io_13_q_reorder = uRegState_13_io_q_reorder; 
  wire [4:0] uRegState_io_12_q_reorder = uRegState_12_io_q_reorder; 
  wire [4:0] uRegState_io_11_q_reorder = uRegState_11_io_q_reorder; 
  wire [4:0] uRegState_io_10_q_reorder = uRegState_10_io_q_reorder; 
  wire [4:0] uRegState_io_9_q_reorder = uRegState_9_io_q_reorder; 
  wire [4:0] uRegState_io_8_q_reorder = uRegState_8_io_q_reorder; 
  wire [4:0] uRegState_io_7_q_reorder = uRegState_7_io_q_reorder; 
  wire [4:0] uRegState_io_6_q_reorder = uRegState_6_io_q_reorder; 
  wire [4:0] uRegState_io_5_q_reorder = uRegState_5_io_q_reorder; 
  wire [4:0] uRegState_io_4_q_reorder = uRegState_4_io_q_reorder; 
  wire [4:0] uRegState_io_3_q_reorder = uRegState_3_io_q_reorder; 
  wire [4:0] uRegState_io_2_q_reorder = uRegState_2_io_q_reorder; 
  wire [4:0] uRegState_io_1_q_reorder = uRegState_1_io_q_reorder; 
  wire [4:0] uRegState_io_0_q_reorder = uRegState_0_io_q_reorder; 
  wire [4:0] _GEN_255 = 5'h1 == decoder_if_rt_idx ? uRegState_io_1_q_reorder : uRegState_io_0_q_reorder; 
  wire [4:0] _GEN_256 = 5'h2 == decoder_if_rt_idx ? uRegState_io_2_q_reorder : _GEN_255; 
  wire [4:0] _GEN_257 = 5'h3 == decoder_if_rt_idx ? uRegState_io_3_q_reorder : _GEN_256; 
  wire [4:0] _GEN_258 = 5'h4 == decoder_if_rt_idx ? uRegState_io_4_q_reorder : _GEN_257; 
  wire [4:0] _GEN_259 = 5'h5 == decoder_if_rt_idx ? uRegState_io_5_q_reorder : _GEN_258; 
  wire [4:0] _GEN_260 = 5'h6 == decoder_if_rt_idx ? uRegState_io_6_q_reorder : _GEN_259; 
  wire [4:0] _GEN_261 = 5'h7 == decoder_if_rt_idx ? uRegState_io_7_q_reorder : _GEN_260; 
  wire [4:0] _GEN_262 = 5'h8 == decoder_if_rt_idx ? uRegState_io_8_q_reorder : _GEN_261; 
  wire [4:0] _GEN_263 = 5'h9 == decoder_if_rt_idx ? uRegState_io_9_q_reorder : _GEN_262; 
  wire [4:0] _GEN_264 = 5'ha == decoder_if_rt_idx ? uRegState_io_10_q_reorder : _GEN_263; 
  wire [4:0] _GEN_265 = 5'hb == decoder_if_rt_idx ? uRegState_io_11_q_reorder : _GEN_264; 
  wire [4:0] _GEN_266 = 5'hc == decoder_if_rt_idx ? uRegState_io_12_q_reorder : _GEN_265; 
  wire [4:0] _GEN_267 = 5'hd == decoder_if_rt_idx ? uRegState_io_13_q_reorder : _GEN_266; 
  wire [4:0] _GEN_268 = 5'he == decoder_if_rt_idx ? uRegState_io_14_q_reorder : _GEN_267; 
  wire [4:0] _GEN_269 = 5'hf == decoder_if_rt_idx ? uRegState_io_15_q_reorder : _GEN_268; 
  wire [4:0] _GEN_270 = 5'h10 == decoder_if_rt_idx ? uRegState_io_16_q_reorder : _GEN_269; 
  wire [4:0] _GEN_271 = 5'h11 == decoder_if_rt_idx ? uRegState_io_17_q_reorder : _GEN_270; 
  wire [4:0] _GEN_272 = 5'h12 == decoder_if_rt_idx ? uRegState_io_18_q_reorder : _GEN_271; 
  wire [4:0] _GEN_273 = 5'h13 == decoder_if_rt_idx ? uRegState_io_19_q_reorder : _GEN_272; 
  wire [4:0] _GEN_274 = 5'h14 == decoder_if_rt_idx ? uRegState_io_20_q_reorder : _GEN_273; 
  wire [4:0] _GEN_275 = 5'h15 == decoder_if_rt_idx ? uRegState_io_21_q_reorder : _GEN_274; 
  wire [4:0] _GEN_276 = 5'h16 == decoder_if_rt_idx ? uRegState_io_22_q_reorder : _GEN_275; 
  wire [4:0] _GEN_277 = 5'h17 == decoder_if_rt_idx ? uRegState_io_23_q_reorder : _GEN_276; 
  wire [4:0] _GEN_278 = 5'h18 == decoder_if_rt_idx ? uRegState_io_24_q_reorder : _GEN_277; 
  wire [4:0] _GEN_279 = 5'h19 == decoder_if_rt_idx ? uRegState_io_25_q_reorder : _GEN_278; 
  wire [4:0] _GEN_280 = 5'h1a == decoder_if_rt_idx ? uRegState_io_26_q_reorder : _GEN_279; 
  wire [4:0] _GEN_281 = 5'h1b == decoder_if_rt_idx ? uRegState_io_27_q_reorder : _GEN_280; 
  wire [4:0] _GEN_282 = 5'h1c == decoder_if_rt_idx ? uRegState_io_28_q_reorder : _GEN_281; 
  wire [4:0] _GEN_283 = 5'h1d == decoder_if_rt_idx ? uRegState_io_29_q_reorder : _GEN_282; 
  wire [4:0] _GEN_284 = 5'h1e == decoder_if_rt_idx ? uRegState_io_30_q_reorder : _GEN_283; 
  wire [4:0] _GEN_285 = 5'h1f == decoder_if_rt_idx ? uRegState_io_31_q_reorder : _GEN_284; 
  wire  _GEN_338 = 5'h1 == _GEN_285 ? uROB_io_queue_data_split_1_rob_ready : uROB_io_queue_data_split_0_rob_ready; 
  wire  _GEN_339 = 5'h2 == _GEN_285 ? uROB_io_queue_data_split_2_rob_ready : _GEN_338; 
  wire  _GEN_340 = 5'h3 == _GEN_285 ? uROB_io_queue_data_split_3_rob_ready : _GEN_339; 
  wire  _GEN_341 = 5'h4 == _GEN_285 ? uROB_io_queue_data_split_4_rob_ready : _GEN_340; 
  wire  _GEN_342 = 5'h5 == _GEN_285 ? uROB_io_queue_data_split_5_rob_ready : _GEN_341; 
  wire  _GEN_343 = 5'h6 == _GEN_285 ? uROB_io_queue_data_split_6_rob_ready : _GEN_342; 
  wire  _GEN_344 = 5'h7 == _GEN_285 ? uROB_io_queue_data_split_7_rob_ready : _GEN_343; 
  wire  _GEN_345 = 5'h8 == _GEN_285 ? uROB_io_queue_data_split_8_rob_ready : _GEN_344; 
  wire  _GEN_346 = 5'h9 == _GEN_285 ? uROB_io_queue_data_split_9_rob_ready : _GEN_345; 
  wire  _GEN_347 = 5'ha == _GEN_285 ? uROB_io_queue_data_split_10_rob_ready : _GEN_346; 
  wire  _GEN_348 = 5'hb == _GEN_285 ? uROB_io_queue_data_split_11_rob_ready : _GEN_347; 
  wire  _GEN_349 = 5'hc == _GEN_285 ? uROB_io_queue_data_split_12_rob_ready : _GEN_348; 
  wire  _GEN_350 = 5'hd == _GEN_285 ? uROB_io_queue_data_split_13_rob_ready : _GEN_349; 
  wire  _GEN_351 = 5'he == _GEN_285 ? uROB_io_queue_data_split_14_rob_ready : _GEN_350; 
  wire  _GEN_352 = 5'hf == _GEN_285 ? uROB_io_queue_data_split_15_rob_ready : _GEN_351; 
  wire  rob_h_rx_1_rob_ready = 5'h10 == _GEN_285 ? uROB_io_queue_data_split_16_rob_ready : _GEN_352; 
  wire [31:0] _GEN_321 = 5'h1 == _GEN_285 ? uROB_io_queue_data_split_1_rob_value : uROB_io_queue_data_split_0_rob_value; 
  wire [31:0] _GEN_322 = 5'h2 == _GEN_285 ? uROB_io_queue_data_split_2_rob_value : _GEN_321; 
  wire [31:0] _GEN_323 = 5'h3 == _GEN_285 ? uROB_io_queue_data_split_3_rob_value : _GEN_322; 
  wire [31:0] _GEN_324 = 5'h4 == _GEN_285 ? uROB_io_queue_data_split_4_rob_value : _GEN_323; 
  wire [31:0] _GEN_325 = 5'h5 == _GEN_285 ? uROB_io_queue_data_split_5_rob_value : _GEN_324; 
  wire [31:0] _GEN_326 = 5'h6 == _GEN_285 ? uROB_io_queue_data_split_6_rob_value : _GEN_325; 
  wire [31:0] _GEN_327 = 5'h7 == _GEN_285 ? uROB_io_queue_data_split_7_rob_value : _GEN_326; 
  wire [31:0] _GEN_328 = 5'h8 == _GEN_285 ? uROB_io_queue_data_split_8_rob_value : _GEN_327; 
  wire [31:0] _GEN_329 = 5'h9 == _GEN_285 ? uROB_io_queue_data_split_9_rob_value : _GEN_328; 
  wire [31:0] _GEN_330 = 5'ha == _GEN_285 ? uROB_io_queue_data_split_10_rob_value : _GEN_329; 
  wire [31:0] _GEN_331 = 5'hb == _GEN_285 ? uROB_io_queue_data_split_11_rob_value : _GEN_330; 
  wire [31:0] _GEN_332 = 5'hc == _GEN_285 ? uROB_io_queue_data_split_12_rob_value : _GEN_331; 
  wire [31:0] _GEN_333 = 5'hd == _GEN_285 ? uROB_io_queue_data_split_13_rob_value : _GEN_332; 
  wire [31:0] _GEN_334 = 5'he == _GEN_285 ? uROB_io_queue_data_split_14_rob_value : _GEN_333; 
  wire [31:0] _GEN_335 = 5'hf == _GEN_285 ? uROB_io_queue_data_split_15_rob_value : _GEN_334; 
  wire [31:0] rob_h_rx_1_rob_value = 5'h10 == _GEN_285 ? uROB_io_queue_data_split_16_rob_value : _GEN_335; 
  wire  _T_362 = uCDB_io_cdb_dest == _GEN_285; 
  wire  _T_363 = uCDB_io_cdb_valid & _T_362; 
  wire [31:0] _GEN_386 = _T_363 ? uCDB_io_cdb_result : 32'h0; 
  wire [31:0] _GEN_388 = rob_h_rx_1_rob_ready ? rob_h_rx_1_rob_value : _GEN_386; 
  wire [31:0] uRegFile_io_31_q = uRegFile_31_io_q; 
  wire [31:0] uRegFile_io_30_q = uRegFile_30_io_q; 
  wire [31:0] uRegFile_io_29_q = uRegFile_29_io_q; 
  wire [31:0] uRegFile_io_28_q = uRegFile_28_io_q; 
  wire [31:0] uRegFile_io_27_q = uRegFile_27_io_q; 
  wire [31:0] uRegFile_io_26_q = uRegFile_26_io_q; 
  wire [31:0] uRegFile_io_25_q = uRegFile_25_io_q; 
  wire [31:0] uRegFile_io_24_q = uRegFile_24_io_q; 
  wire [31:0] uRegFile_io_23_q = uRegFile_23_io_q; 
  wire [31:0] uRegFile_io_22_q = uRegFile_22_io_q; 
  wire [31:0] uRegFile_io_21_q = uRegFile_21_io_q; 
  wire [31:0] uRegFile_io_20_q = uRegFile_20_io_q; 
  wire [31:0] uRegFile_io_19_q = uRegFile_19_io_q; 
  wire [31:0] uRegFile_io_18_q = uRegFile_18_io_q; 
  wire [31:0] uRegFile_io_17_q = uRegFile_17_io_q; 
  wire [31:0] uRegFile_io_16_q = uRegFile_16_io_q; 
  wire [31:0] uRegFile_io_15_q = uRegFile_15_io_q; 
  wire [31:0] uRegFile_io_14_q = uRegFile_14_io_q; 
  wire [31:0] uRegFile_io_13_q = uRegFile_13_io_q; 
  wire [31:0] uRegFile_io_12_q = uRegFile_12_io_q; 
  wire [31:0] uRegFile_io_11_q = uRegFile_11_io_q; 
  wire [31:0] uRegFile_io_10_q = uRegFile_10_io_q; 
  wire [31:0] uRegFile_io_9_q = uRegFile_9_io_q; 
  wire [31:0] uRegFile_io_8_q = uRegFile_8_io_q; 
  wire [31:0] uRegFile_io_7_q = uRegFile_7_io_q; 
  wire [31:0] uRegFile_io_6_q = uRegFile_6_io_q; 
  wire [31:0] uRegFile_io_5_q = uRegFile_5_io_q; 
  wire [31:0] uRegFile_io_4_q = uRegFile_4_io_q; 
  wire [31:0] uRegFile_io_3_q = uRegFile_3_io_q; 
  wire [31:0] uRegFile_io_2_q = uRegFile_2_io_q; 
  wire [31:0] uRegFile_io_1_q = uRegFile_1_io_q; 
  wire [31:0] uRegFile_io_0_q = uRegFile_0_io_q; 
  wire [31:0] _GEN_391 = 5'h1 == decoder_if_rt_idx ? uRegFile_io_1_q : uRegFile_io_0_q; 
  wire [31:0] _GEN_392 = 5'h2 == decoder_if_rt_idx ? uRegFile_io_2_q : _GEN_391; 
  wire [31:0] _GEN_393 = 5'h3 == decoder_if_rt_idx ? uRegFile_io_3_q : _GEN_392; 
  wire [31:0] _GEN_394 = 5'h4 == decoder_if_rt_idx ? uRegFile_io_4_q : _GEN_393; 
  wire [31:0] _GEN_395 = 5'h5 == decoder_if_rt_idx ? uRegFile_io_5_q : _GEN_394; 
  wire [31:0] _GEN_396 = 5'h6 == decoder_if_rt_idx ? uRegFile_io_6_q : _GEN_395; 
  wire [31:0] _GEN_397 = 5'h7 == decoder_if_rt_idx ? uRegFile_io_7_q : _GEN_396; 
  wire [31:0] _GEN_398 = 5'h8 == decoder_if_rt_idx ? uRegFile_io_8_q : _GEN_397; 
  wire [31:0] _GEN_399 = 5'h9 == decoder_if_rt_idx ? uRegFile_io_9_q : _GEN_398; 
  wire [31:0] _GEN_400 = 5'ha == decoder_if_rt_idx ? uRegFile_io_10_q : _GEN_399; 
  wire [31:0] _GEN_401 = 5'hb == decoder_if_rt_idx ? uRegFile_io_11_q : _GEN_400; 
  wire [31:0] _GEN_402 = 5'hc == decoder_if_rt_idx ? uRegFile_io_12_q : _GEN_401; 
  wire [31:0] _GEN_403 = 5'hd == decoder_if_rt_idx ? uRegFile_io_13_q : _GEN_402; 
  wire [31:0] _GEN_404 = 5'he == decoder_if_rt_idx ? uRegFile_io_14_q : _GEN_403; 
  wire [31:0] _GEN_405 = 5'hf == decoder_if_rt_idx ? uRegFile_io_15_q : _GEN_404; 
  wire [31:0] _GEN_406 = 5'h10 == decoder_if_rt_idx ? uRegFile_io_16_q : _GEN_405; 
  wire [31:0] _GEN_407 = 5'h11 == decoder_if_rt_idx ? uRegFile_io_17_q : _GEN_406; 
  wire [31:0] _GEN_408 = 5'h12 == decoder_if_rt_idx ? uRegFile_io_18_q : _GEN_407; 
  wire [31:0] _GEN_409 = 5'h13 == decoder_if_rt_idx ? uRegFile_io_19_q : _GEN_408; 
  wire [31:0] _GEN_410 = 5'h14 == decoder_if_rt_idx ? uRegFile_io_20_q : _GEN_409; 
  wire [31:0] _GEN_411 = 5'h15 == decoder_if_rt_idx ? uRegFile_io_21_q : _GEN_410; 
  wire [31:0] _GEN_412 = 5'h16 == decoder_if_rt_idx ? uRegFile_io_22_q : _GEN_411; 
  wire [31:0] _GEN_413 = 5'h17 == decoder_if_rt_idx ? uRegFile_io_23_q : _GEN_412; 
  wire [31:0] _GEN_414 = 5'h18 == decoder_if_rt_idx ? uRegFile_io_24_q : _GEN_413; 
  wire [31:0] _GEN_415 = 5'h19 == decoder_if_rt_idx ? uRegFile_io_25_q : _GEN_414; 
  wire [31:0] _GEN_416 = 5'h1a == decoder_if_rt_idx ? uRegFile_io_26_q : _GEN_415; 
  wire [31:0] _GEN_417 = 5'h1b == decoder_if_rt_idx ? uRegFile_io_27_q : _GEN_416; 
  wire [31:0] _GEN_418 = 5'h1c == decoder_if_rt_idx ? uRegFile_io_28_q : _GEN_417; 
  wire [31:0] _GEN_419 = 5'h1d == decoder_if_rt_idx ? uRegFile_io_29_q : _GEN_418; 
  wire [31:0] _GEN_420 = 5'h1e == decoder_if_rt_idx ? uRegFile_io_30_q : _GEN_419; 
  wire [31:0] _GEN_421 = 5'h1f == decoder_if_rt_idx ? uRegFile_io_31_q : _GEN_420; 
  wire [31:0] _GEN_422 = _GEN_385 ? _GEN_388 : _GEN_421; 
  wire [31:0] _GEN_424 = decoder_if_exe_op_jr ? decoder_if_pc_out : decoder_if_imm; 
  wire [31:0] _GEN_425 = decoder_if_rt_idx_valid ? _GEN_422 : _GEN_424; 
  wire [31:0] _GEN_499 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_425 : 32'h0; 
  wire [31:0] _GEN_913 = _T_352 ? _GEN_422 : 32'h0; 
  wire [31:0] _GEN_2334 = branch_inst_r_io_d ? _GEN_913 : 32'h0; 
  wire [31:0] _GEN_2424 = integer_inst_r_io_d ? _GEN_499 : _GEN_2334; 
  wire [31:0] uIntergerRS_io_enq_data_vk = decoder_if_inst_valid ? _GEN_2424 : 32'h0; 
  wire  _GEN_2329 = branch_inst_r_io_d & _T_352; 
  wire  _GEN_2419 = integer_inst_r_io_d ? _T_352 : _GEN_2329; 
  wire  uIntergerRS_io_enq_data_busy = decoder_if_inst_valid & _GEN_2419; 
  wire  _GEN_185 = 5'h1 == decoder_if_rs_idx ? uRegState_io_1_q_busy : uRegState_io_0_q_busy; 
  wire  _GEN_186 = 5'h2 == decoder_if_rs_idx ? uRegState_io_2_q_busy : _GEN_185; 
  wire  _GEN_187 = 5'h3 == decoder_if_rs_idx ? uRegState_io_3_q_busy : _GEN_186; 
  wire  _GEN_188 = 5'h4 == decoder_if_rs_idx ? uRegState_io_4_q_busy : _GEN_187; 
  wire  _GEN_189 = 5'h5 == decoder_if_rs_idx ? uRegState_io_5_q_busy : _GEN_188; 
  wire  _GEN_190 = 5'h6 == decoder_if_rs_idx ? uRegState_io_6_q_busy : _GEN_189; 
  wire  _GEN_191 = 5'h7 == decoder_if_rs_idx ? uRegState_io_7_q_busy : _GEN_190; 
  wire  _GEN_192 = 5'h8 == decoder_if_rs_idx ? uRegState_io_8_q_busy : _GEN_191; 
  wire  _GEN_193 = 5'h9 == decoder_if_rs_idx ? uRegState_io_9_q_busy : _GEN_192; 
  wire  _GEN_194 = 5'ha == decoder_if_rs_idx ? uRegState_io_10_q_busy : _GEN_193; 
  wire  _GEN_195 = 5'hb == decoder_if_rs_idx ? uRegState_io_11_q_busy : _GEN_194; 
  wire  _GEN_196 = 5'hc == decoder_if_rs_idx ? uRegState_io_12_q_busy : _GEN_195; 
  wire  _GEN_197 = 5'hd == decoder_if_rs_idx ? uRegState_io_13_q_busy : _GEN_196; 
  wire  _GEN_198 = 5'he == decoder_if_rs_idx ? uRegState_io_14_q_busy : _GEN_197; 
  wire  _GEN_199 = 5'hf == decoder_if_rs_idx ? uRegState_io_15_q_busy : _GEN_198; 
  wire  _GEN_200 = 5'h10 == decoder_if_rs_idx ? uRegState_io_16_q_busy : _GEN_199; 
  wire  _GEN_201 = 5'h11 == decoder_if_rs_idx ? uRegState_io_17_q_busy : _GEN_200; 
  wire  _GEN_202 = 5'h12 == decoder_if_rs_idx ? uRegState_io_18_q_busy : _GEN_201; 
  wire  _GEN_203 = 5'h13 == decoder_if_rs_idx ? uRegState_io_19_q_busy : _GEN_202; 
  wire  _GEN_204 = 5'h14 == decoder_if_rs_idx ? uRegState_io_20_q_busy : _GEN_203; 
  wire  _GEN_205 = 5'h15 == decoder_if_rs_idx ? uRegState_io_21_q_busy : _GEN_204; 
  wire  _GEN_206 = 5'h16 == decoder_if_rs_idx ? uRegState_io_22_q_busy : _GEN_205; 
  wire  _GEN_207 = 5'h17 == decoder_if_rs_idx ? uRegState_io_23_q_busy : _GEN_206; 
  wire  _GEN_208 = 5'h18 == decoder_if_rs_idx ? uRegState_io_24_q_busy : _GEN_207; 
  wire  _GEN_209 = 5'h19 == decoder_if_rs_idx ? uRegState_io_25_q_busy : _GEN_208; 
  wire  _GEN_210 = 5'h1a == decoder_if_rs_idx ? uRegState_io_26_q_busy : _GEN_209; 
  wire  _GEN_211 = 5'h1b == decoder_if_rs_idx ? uRegState_io_27_q_busy : _GEN_210; 
  wire  _GEN_212 = 5'h1c == decoder_if_rs_idx ? uRegState_io_28_q_busy : _GEN_211; 
  wire  _GEN_213 = 5'h1d == decoder_if_rs_idx ? uRegState_io_29_q_busy : _GEN_212; 
  wire  _GEN_214 = 5'h1e == decoder_if_rs_idx ? uRegState_io_30_q_busy : _GEN_213; 
  wire  _GEN_215 = 5'h1f == decoder_if_rs_idx ? uRegState_io_31_q_busy : _GEN_214; 
  wire [4:0] _GEN_85 = 5'h1 == decoder_if_rs_idx ? uRegState_io_1_q_reorder : uRegState_io_0_q_reorder; 
  wire [4:0] _GEN_86 = 5'h2 == decoder_if_rs_idx ? uRegState_io_2_q_reorder : _GEN_85; 
  wire [4:0] _GEN_87 = 5'h3 == decoder_if_rs_idx ? uRegState_io_3_q_reorder : _GEN_86; 
  wire [4:0] _GEN_88 = 5'h4 == decoder_if_rs_idx ? uRegState_io_4_q_reorder : _GEN_87; 
  wire [4:0] _GEN_89 = 5'h5 == decoder_if_rs_idx ? uRegState_io_5_q_reorder : _GEN_88; 
  wire [4:0] _GEN_90 = 5'h6 == decoder_if_rs_idx ? uRegState_io_6_q_reorder : _GEN_89; 
  wire [4:0] _GEN_91 = 5'h7 == decoder_if_rs_idx ? uRegState_io_7_q_reorder : _GEN_90; 
  wire [4:0] _GEN_92 = 5'h8 == decoder_if_rs_idx ? uRegState_io_8_q_reorder : _GEN_91; 
  wire [4:0] _GEN_93 = 5'h9 == decoder_if_rs_idx ? uRegState_io_9_q_reorder : _GEN_92; 
  wire [4:0] _GEN_94 = 5'ha == decoder_if_rs_idx ? uRegState_io_10_q_reorder : _GEN_93; 
  wire [4:0] _GEN_95 = 5'hb == decoder_if_rs_idx ? uRegState_io_11_q_reorder : _GEN_94; 
  wire [4:0] _GEN_96 = 5'hc == decoder_if_rs_idx ? uRegState_io_12_q_reorder : _GEN_95; 
  wire [4:0] _GEN_97 = 5'hd == decoder_if_rs_idx ? uRegState_io_13_q_reorder : _GEN_96; 
  wire [4:0] _GEN_98 = 5'he == decoder_if_rs_idx ? uRegState_io_14_q_reorder : _GEN_97; 
  wire [4:0] _GEN_99 = 5'hf == decoder_if_rs_idx ? uRegState_io_15_q_reorder : _GEN_98; 
  wire [4:0] _GEN_100 = 5'h10 == decoder_if_rs_idx ? uRegState_io_16_q_reorder : _GEN_99; 
  wire [4:0] _GEN_101 = 5'h11 == decoder_if_rs_idx ? uRegState_io_17_q_reorder : _GEN_100; 
  wire [4:0] _GEN_102 = 5'h12 == decoder_if_rs_idx ? uRegState_io_18_q_reorder : _GEN_101; 
  wire [4:0] _GEN_103 = 5'h13 == decoder_if_rs_idx ? uRegState_io_19_q_reorder : _GEN_102; 
  wire [4:0] _GEN_104 = 5'h14 == decoder_if_rs_idx ? uRegState_io_20_q_reorder : _GEN_103; 
  wire [4:0] _GEN_105 = 5'h15 == decoder_if_rs_idx ? uRegState_io_21_q_reorder : _GEN_104; 
  wire [4:0] _GEN_106 = 5'h16 == decoder_if_rs_idx ? uRegState_io_22_q_reorder : _GEN_105; 
  wire [4:0] _GEN_107 = 5'h17 == decoder_if_rs_idx ? uRegState_io_23_q_reorder : _GEN_106; 
  wire [4:0] _GEN_108 = 5'h18 == decoder_if_rs_idx ? uRegState_io_24_q_reorder : _GEN_107; 
  wire [4:0] _GEN_109 = 5'h19 == decoder_if_rs_idx ? uRegState_io_25_q_reorder : _GEN_108; 
  wire [4:0] _GEN_110 = 5'h1a == decoder_if_rs_idx ? uRegState_io_26_q_reorder : _GEN_109; 
  wire [4:0] _GEN_111 = 5'h1b == decoder_if_rs_idx ? uRegState_io_27_q_reorder : _GEN_110; 
  wire [4:0] _GEN_112 = 5'h1c == decoder_if_rs_idx ? uRegState_io_28_q_reorder : _GEN_111; 
  wire [4:0] _GEN_113 = 5'h1d == decoder_if_rs_idx ? uRegState_io_29_q_reorder : _GEN_112; 
  wire [4:0] _GEN_114 = 5'h1e == decoder_if_rs_idx ? uRegState_io_30_q_reorder : _GEN_113; 
  wire [4:0] _GEN_115 = 5'h1f == decoder_if_rs_idx ? uRegState_io_31_q_reorder : _GEN_114; 
  wire  _GEN_168 = 5'h1 == _GEN_115 ? uROB_io_queue_data_split_1_rob_ready : uROB_io_queue_data_split_0_rob_ready; 
  wire  _GEN_169 = 5'h2 == _GEN_115 ? uROB_io_queue_data_split_2_rob_ready : _GEN_168; 
  wire  _GEN_170 = 5'h3 == _GEN_115 ? uROB_io_queue_data_split_3_rob_ready : _GEN_169; 
  wire  _GEN_171 = 5'h4 == _GEN_115 ? uROB_io_queue_data_split_4_rob_ready : _GEN_170; 
  wire  _GEN_172 = 5'h5 == _GEN_115 ? uROB_io_queue_data_split_5_rob_ready : _GEN_171; 
  wire  _GEN_173 = 5'h6 == _GEN_115 ? uROB_io_queue_data_split_6_rob_ready : _GEN_172; 
  wire  _GEN_174 = 5'h7 == _GEN_115 ? uROB_io_queue_data_split_7_rob_ready : _GEN_173; 
  wire  _GEN_175 = 5'h8 == _GEN_115 ? uROB_io_queue_data_split_8_rob_ready : _GEN_174; 
  wire  _GEN_176 = 5'h9 == _GEN_115 ? uROB_io_queue_data_split_9_rob_ready : _GEN_175; 
  wire  _GEN_177 = 5'ha == _GEN_115 ? uROB_io_queue_data_split_10_rob_ready : _GEN_176; 
  wire  _GEN_178 = 5'hb == _GEN_115 ? uROB_io_queue_data_split_11_rob_ready : _GEN_177; 
  wire  _GEN_179 = 5'hc == _GEN_115 ? uROB_io_queue_data_split_12_rob_ready : _GEN_178; 
  wire  _GEN_180 = 5'hd == _GEN_115 ? uROB_io_queue_data_split_13_rob_ready : _GEN_179; 
  wire  _GEN_181 = 5'he == _GEN_115 ? uROB_io_queue_data_split_14_rob_ready : _GEN_180; 
  wire  _GEN_182 = 5'hf == _GEN_115 ? uROB_io_queue_data_split_15_rob_ready : _GEN_181; 
  wire  rob_h_rx_rob_ready = 5'h10 == _GEN_115 ? uROB_io_queue_data_split_16_rob_ready : _GEN_182; 
  wire [31:0] _GEN_151 = 5'h1 == _GEN_115 ? uROB_io_queue_data_split_1_rob_value : uROB_io_queue_data_split_0_rob_value; 
  wire [31:0] _GEN_152 = 5'h2 == _GEN_115 ? uROB_io_queue_data_split_2_rob_value : _GEN_151; 
  wire [31:0] _GEN_153 = 5'h3 == _GEN_115 ? uROB_io_queue_data_split_3_rob_value : _GEN_152; 
  wire [31:0] _GEN_154 = 5'h4 == _GEN_115 ? uROB_io_queue_data_split_4_rob_value : _GEN_153; 
  wire [31:0] _GEN_155 = 5'h5 == _GEN_115 ? uROB_io_queue_data_split_5_rob_value : _GEN_154; 
  wire [31:0] _GEN_156 = 5'h6 == _GEN_115 ? uROB_io_queue_data_split_6_rob_value : _GEN_155; 
  wire [31:0] _GEN_157 = 5'h7 == _GEN_115 ? uROB_io_queue_data_split_7_rob_value : _GEN_156; 
  wire [31:0] _GEN_158 = 5'h8 == _GEN_115 ? uROB_io_queue_data_split_8_rob_value : _GEN_157; 
  wire [31:0] _GEN_159 = 5'h9 == _GEN_115 ? uROB_io_queue_data_split_9_rob_value : _GEN_158; 
  wire [31:0] _GEN_160 = 5'ha == _GEN_115 ? uROB_io_queue_data_split_10_rob_value : _GEN_159; 
  wire [31:0] _GEN_161 = 5'hb == _GEN_115 ? uROB_io_queue_data_split_11_rob_value : _GEN_160; 
  wire [31:0] _GEN_162 = 5'hc == _GEN_115 ? uROB_io_queue_data_split_12_rob_value : _GEN_161; 
  wire [31:0] _GEN_163 = 5'hd == _GEN_115 ? uROB_io_queue_data_split_13_rob_value : _GEN_162; 
  wire [31:0] _GEN_164 = 5'he == _GEN_115 ? uROB_io_queue_data_split_14_rob_value : _GEN_163; 
  wire [31:0] _GEN_165 = 5'hf == _GEN_115 ? uROB_io_queue_data_split_15_rob_value : _GEN_164; 
  wire [31:0] rob_h_rx_rob_value = 5'h10 == _GEN_115 ? uROB_io_queue_data_split_16_rob_value : _GEN_165; 
  wire  _T_356 = uCDB_io_cdb_dest == _GEN_115; 
  wire  _T_357 = uCDB_io_cdb_valid & _T_356; 
  wire [31:0] _GEN_216 = _T_357 ? uCDB_io_cdb_result : 32'h0; 
  wire [31:0] _GEN_218 = rob_h_rx_rob_ready ? rob_h_rx_rob_value : _GEN_216; 
  wire [31:0] _GEN_221 = 5'h1 == decoder_if_rs_idx ? uRegFile_io_1_q : uRegFile_io_0_q; 
  wire [31:0] _GEN_222 = 5'h2 == decoder_if_rs_idx ? uRegFile_io_2_q : _GEN_221; 
  wire [31:0] _GEN_223 = 5'h3 == decoder_if_rs_idx ? uRegFile_io_3_q : _GEN_222; 
  wire [31:0] _GEN_224 = 5'h4 == decoder_if_rs_idx ? uRegFile_io_4_q : _GEN_223; 
  wire [31:0] _GEN_225 = 5'h5 == decoder_if_rs_idx ? uRegFile_io_5_q : _GEN_224; 
  wire [31:0] _GEN_226 = 5'h6 == decoder_if_rs_idx ? uRegFile_io_6_q : _GEN_225; 
  wire [31:0] _GEN_227 = 5'h7 == decoder_if_rs_idx ? uRegFile_io_7_q : _GEN_226; 
  wire [31:0] _GEN_228 = 5'h8 == decoder_if_rs_idx ? uRegFile_io_8_q : _GEN_227; 
  wire [31:0] _GEN_229 = 5'h9 == decoder_if_rs_idx ? uRegFile_io_9_q : _GEN_228; 
  wire [31:0] _GEN_230 = 5'ha == decoder_if_rs_idx ? uRegFile_io_10_q : _GEN_229; 
  wire [31:0] _GEN_231 = 5'hb == decoder_if_rs_idx ? uRegFile_io_11_q : _GEN_230; 
  wire [31:0] _GEN_232 = 5'hc == decoder_if_rs_idx ? uRegFile_io_12_q : _GEN_231; 
  wire [31:0] _GEN_233 = 5'hd == decoder_if_rs_idx ? uRegFile_io_13_q : _GEN_232; 
  wire [31:0] _GEN_234 = 5'he == decoder_if_rs_idx ? uRegFile_io_14_q : _GEN_233; 
  wire [31:0] _GEN_235 = 5'hf == decoder_if_rs_idx ? uRegFile_io_15_q : _GEN_234; 
  wire [31:0] _GEN_236 = 5'h10 == decoder_if_rs_idx ? uRegFile_io_16_q : _GEN_235; 
  wire [31:0] _GEN_237 = 5'h11 == decoder_if_rs_idx ? uRegFile_io_17_q : _GEN_236; 
  wire [31:0] _GEN_238 = 5'h12 == decoder_if_rs_idx ? uRegFile_io_18_q : _GEN_237; 
  wire [31:0] _GEN_239 = 5'h13 == decoder_if_rs_idx ? uRegFile_io_19_q : _GEN_238; 
  wire [31:0] _GEN_240 = 5'h14 == decoder_if_rs_idx ? uRegFile_io_20_q : _GEN_239; 
  wire [31:0] _GEN_241 = 5'h15 == decoder_if_rs_idx ? uRegFile_io_21_q : _GEN_240; 
  wire [31:0] _GEN_242 = 5'h16 == decoder_if_rs_idx ? uRegFile_io_22_q : _GEN_241; 
  wire [31:0] _GEN_243 = 5'h17 == decoder_if_rs_idx ? uRegFile_io_23_q : _GEN_242; 
  wire [31:0] _GEN_244 = 5'h18 == decoder_if_rs_idx ? uRegFile_io_24_q : _GEN_243; 
  wire [31:0] _GEN_245 = 5'h19 == decoder_if_rs_idx ? uRegFile_io_25_q : _GEN_244; 
  wire [31:0] _GEN_246 = 5'h1a == decoder_if_rs_idx ? uRegFile_io_26_q : _GEN_245; 
  wire [31:0] _GEN_247 = 5'h1b == decoder_if_rs_idx ? uRegFile_io_27_q : _GEN_246; 
  wire [31:0] _GEN_248 = 5'h1c == decoder_if_rs_idx ? uRegFile_io_28_q : _GEN_247; 
  wire [31:0] _GEN_249 = 5'h1d == decoder_if_rs_idx ? uRegFile_io_29_q : _GEN_248; 
  wire [31:0] _GEN_250 = 5'h1e == decoder_if_rs_idx ? uRegFile_io_30_q : _GEN_249; 
  wire [31:0] _GEN_251 = 5'h1f == decoder_if_rs_idx ? uRegFile_io_31_q : _GEN_250; 
  wire [31:0] _GEN_252 = _GEN_215 ? _GEN_218 : _GEN_251; 
  wire [31:0] _GEN_497 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_252 : 32'h0; 
  wire [31:0] _GEN_2332 = branch_inst_r_io_d ? _GEN_497 : 32'h0; 
  wire [31:0] _GEN_2422 = integer_inst_r_io_d ? _GEN_497 : _GEN_2332; 
  wire [31:0] uIntergerRS_io_enq_data_vj = decoder_if_inst_valid ? _GEN_2422 : 32'h0; 
  wire [96:0] uIntergerRS_io_enq_data_lo = {32'h0,uIntergerRS_io_enq_data_vj,uIntergerRS_io_enq_data_vk,
    uIntergerRS_io_enq_data_busy}; 
  wire [4:0] _GEN_217 = _T_357 ? 5'h0 : _GEN_115; 
  wire [4:0] _GEN_219 = rob_h_rx_rob_ready ? 5'h0 : _GEN_217; 
  wire [4:0] _GEN_253 = _GEN_215 ? _GEN_219 : 5'h0; 
  wire [4:0] _GEN_498 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_253 : 5'h0; 
  wire [4:0] _GEN_2333 = branch_inst_r_io_d ? _GEN_498 : 5'h0; 
  wire [4:0] _GEN_2423 = integer_inst_r_io_d ? _GEN_498 : _GEN_2333; 
  wire [4:0] uIntergerRS_io_enq_data_qj = decoder_if_inst_valid ? _GEN_2423 : 5'h0; 
  wire [4:0] _GEN_387 = _T_363 ? 5'h0 : _GEN_285; 
  wire [4:0] _GEN_389 = rob_h_rx_1_rob_ready ? 5'h0 : _GEN_387; 
  wire [4:0] _GEN_423 = _GEN_385 ? _GEN_389 : 5'h0; 
  wire [4:0] _GEN_426 = decoder_if_rt_idx_valid ? _GEN_423 : 5'h0; 
  wire [4:0] _GEN_500 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_426 : 5'h0; 
  wire [4:0] _GEN_914 = _T_352 ? _GEN_423 : 5'h0; 
  wire [4:0] _GEN_2335 = branch_inst_r_io_d ? _GEN_914 : 5'h0; 
  wire [4:0] _GEN_2425 = integer_inst_r_io_d ? _GEN_500 : _GEN_2335; 
  wire [4:0] uIntergerRS_io_enq_data_qk = decoder_if_inst_valid ? _GEN_2425 : 5'h0; 
  wire [9:0] uIntergerRS_io_enq_data_op_hi = {decoder_if_exe_op_store,decoder_if_exe_op_load,decoder_if_exe_op_muldivb_s
    ,decoder_if_exe_op_muldiva_s,decoder_if_exe_op_div,decoder_if_exe_op_mul,decoder_if_exe_op_equal,
    decoder_if_exe_op_large,decoder_if_exe_op_less,decoder_if_exe_op_jr}; 
  wire [9:0] uIntergerRS_io_enq_data_op_lo = {decoder_if_exe_op_br,decoder_if_exe_op_sra,decoder_if_exe_op_srl,
    decoder_if_exe_op_sll,decoder_if_exe_op_sub,decoder_if_exe_op_add,decoder_if_exe_op_set,decoder_if_exe_op_xor,
    decoder_if_exe_op_or,decoder_if_exe_op_and}; 
  wire [19:0] _uIntergerRS_io_enq_data_op_T = {uIntergerRS_io_enq_data_op_hi,uIntergerRS_io_enq_data_op_lo}; 
  wire [19:0] _GEN_495 = ~uIntergerRS__io_full & ~uROB__io_full ? _uIntergerRS_io_enq_data_op_T : 20'h0; 
  wire [19:0] _GEN_2330 = branch_inst_r_io_d ? _GEN_495 : 20'h0; 
  wire [19:0] _GEN_2420 = integer_inst_r_io_d ? _GEN_495 : _GEN_2330; 
  wire [19:0] uIntergerRS_io_enq_data_op = decoder_if_inst_valid ? _GEN_2420 : 20'h0; 
  wire [4:0] _GEN_496 = ~uIntergerRS__io_full & ~uROB__io_full ? uROB__io_enq_idx : 5'h0; 
  wire [4:0] _GEN_2331 = branch_inst_r_io_d ? _GEN_496 : 5'h0; 
  wire [4:0] _GEN_2421 = integer_inst_r_io_d ? _GEN_496 : _GEN_2331; 
  wire [4:0] uIntergerRS_io_enq_data_dest = decoder_if_inst_valid ? _GEN_2421 : 5'h0; 
  wire [34:0] uIntergerRS_io_enq_data_hi = {uIntergerRS_io_enq_data_op,uIntergerRS_io_enq_data_dest,
    uIntergerRS_io_enq_data_qj,uIntergerRS_io_enq_data_qk}; 
  wire [19:0] uIntergerRS_io_deq_data_op = uIntergerRS__io_deq_data[131:112]; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_1 = uIntergerRS_io_queue_data_split_1_qj == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_2 = ~uIntergerRS__io_empty & _uIntergerRS_io_deq_cond_vec_1_T_1; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_3 = uIntergerRS_io_queue_data_split_1_qk == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_4 = _uIntergerRS_io_deq_cond_vec_1_T_2 & _uIntergerRS_io_deq_cond_vec_1_T_3; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_6 = _uIntergerRS_io_deq_cond_vec_1_T_4 & uIntergerRS_io_queue_data_split_1_busy
    ; 
  wire  _uIntergerRS_io_deq_cond_vec_1_T_8 = ~uIntBusGetData_st_io_q | uCDB_io_int_ready; 
  wire  uIntergerRS_io_deq_cond_vec_1 = _uIntergerRS_io_deq_cond_vec_1_T_6 & _uIntergerRS_io_deq_cond_vec_1_T_8; 
  wire  _uIntergerRS_io_deq_cond_vec_0_T_1 = uIntergerRS_io_queue_data_split_0_qj == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_0_T_2 = ~uIntergerRS__io_empty & _uIntergerRS_io_deq_cond_vec_0_T_1; 
  wire  _uIntergerRS_io_deq_cond_vec_0_T_3 = uIntergerRS_io_queue_data_split_0_qk == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_0_T_4 = _uIntergerRS_io_deq_cond_vec_0_T_2 & _uIntergerRS_io_deq_cond_vec_0_T_3; 
  wire  _uIntergerRS_io_deq_cond_vec_0_T_6 = _uIntergerRS_io_deq_cond_vec_0_T_4 & uIntergerRS_io_queue_data_split_0_busy
    ; 
  wire  uIntergerRS_io_deq_cond_vec_0 = _uIntergerRS_io_deq_cond_vec_0_T_6 & _uIntergerRS_io_deq_cond_vec_1_T_8; 
  wire [1:0] uIntergerRS_io_deq_cond_lo = {uIntergerRS_io_deq_cond_vec_1,uIntergerRS_io_deq_cond_vec_0}; 
  wire  _uIntergerRS_io_deq_cond_vec_3_T_1 = uIntergerRS_io_queue_data_split_3_qj == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_3_T_2 = ~uIntergerRS__io_empty & _uIntergerRS_io_deq_cond_vec_3_T_1; 
  wire  _uIntergerRS_io_deq_cond_vec_3_T_3 = uIntergerRS_io_queue_data_split_3_qk == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_3_T_4 = _uIntergerRS_io_deq_cond_vec_3_T_2 & _uIntergerRS_io_deq_cond_vec_3_T_3; 
  wire  _uIntergerRS_io_deq_cond_vec_3_T_6 = _uIntergerRS_io_deq_cond_vec_3_T_4 & uIntergerRS_io_queue_data_split_3_busy
    ; 
  wire  uIntergerRS_io_deq_cond_vec_3 = _uIntergerRS_io_deq_cond_vec_3_T_6 & _uIntergerRS_io_deq_cond_vec_1_T_8; 
  wire  _uIntergerRS_io_deq_cond_vec_2_T_1 = uIntergerRS_io_queue_data_split_2_qj == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_2_T_2 = ~uIntergerRS__io_empty & _uIntergerRS_io_deq_cond_vec_2_T_1; 
  wire  _uIntergerRS_io_deq_cond_vec_2_T_3 = uIntergerRS_io_queue_data_split_2_qk == 5'h0; 
  wire  _uIntergerRS_io_deq_cond_vec_2_T_4 = _uIntergerRS_io_deq_cond_vec_2_T_2 & _uIntergerRS_io_deq_cond_vec_2_T_3; 
  wire  _uIntergerRS_io_deq_cond_vec_2_T_6 = _uIntergerRS_io_deq_cond_vec_2_T_4 & uIntergerRS_io_queue_data_split_2_busy
    ; 
  wire  uIntergerRS_io_deq_cond_vec_2 = _uIntergerRS_io_deq_cond_vec_2_T_6 & _uIntergerRS_io_deq_cond_vec_1_T_8; 
  wire [1:0] uIntergerRS_io_deq_cond_hi = {uIntergerRS_io_deq_cond_vec_3,uIntergerRS_io_deq_cond_vec_2}; 
  wire  _T_529 = uCDB_io_cdb_valid; 
  wire  _T_530 = uIntergerRS_io_queue_data_split_1_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qj_entry_1 = uCDB_io_cdb_valid & _T_530; 
  wire  _T_532 = uIntergerRS_io_queue_data_split_1_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qk_entry_1 = uCDB_io_cdb_valid & _T_532; 
  wire  _T_534 = need2_update_uIntegerRS_Qj_entry_1 | need2_update_uIntegerRS_Qk_entry_1; 
  wire  uIntergerRS_io_update_entry_1 = uCDB_io_cdb_valid & _T_534; 
  wire  _T_521 = uIntergerRS_io_queue_data_split_0_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qj_entry_0 = uCDB_io_cdb_valid & _T_521; 
  wire  _T_523 = uIntergerRS_io_queue_data_split_0_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qk_entry_0 = uCDB_io_cdb_valid & _T_523; 
  wire  _T_525 = need2_update_uIntegerRS_Qj_entry_0 | need2_update_uIntegerRS_Qk_entry_0; 
  wire  uIntergerRS_io_update_entry_0 = uCDB_io_cdb_valid & _T_525; 
  wire [1:0] uIntergerRS_io_update_entry_lo = {uIntergerRS_io_update_entry_1,uIntergerRS_io_update_entry_0}; 
  wire  _T_548 = uIntergerRS_io_queue_data_split_3_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qj_entry_3 = uCDB_io_cdb_valid & _T_548; 
  wire  _T_550 = uIntergerRS_io_queue_data_split_3_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qk_entry_3 = uCDB_io_cdb_valid & _T_550; 
  wire  _T_552 = need2_update_uIntegerRS_Qj_entry_3 | need2_update_uIntegerRS_Qk_entry_3; 
  wire  uIntergerRS_io_update_entry_3 = uCDB_io_cdb_valid & _T_552; 
  wire  _T_539 = uIntergerRS_io_queue_data_split_2_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qj_entry_2 = uCDB_io_cdb_valid & _T_539; 
  wire  _T_541 = uIntergerRS_io_queue_data_split_2_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uIntegerRS_Qk_entry_2 = uCDB_io_cdb_valid & _T_541; 
  wire  _T_543 = need2_update_uIntegerRS_Qj_entry_2 | need2_update_uIntegerRS_Qk_entry_2; 
  wire  uIntergerRS_io_update_entry_2 = uCDB_io_cdb_valid & _T_543; 
  wire [1:0] uIntergerRS_io_update_entry_hi = {uIntergerRS_io_update_entry_3,uIntergerRS_io_update_entry_2}; 
  wire [31:0] _GEN_2764 = need2_update_uIntegerRS_Qk_entry_0 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_0_vk
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_0_vk = uCDB_io_cdb_valid ? _GEN_2764 :
    uIntergerRS_io_queue_data_split_0_vk; 
  wire [31:0] _GEN_2762 = need2_update_uIntegerRS_Qj_entry_0 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_0_vj
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_0_vj = uCDB_io_cdb_valid ? _GEN_2762 :
    uIntergerRS_io_queue_data_split_0_vj; 
  wire [4:0] _GEN_2761 = need2_update_uIntegerRS_Qj_entry_0 ? 5'h0 : uIntergerRS_io_queue_data_split_0_qj; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_0_qj = uCDB_io_cdb_valid ? _GEN_2761 :
    uIntergerRS_io_queue_data_split_0_qj; 
  wire [4:0] _GEN_2763 = need2_update_uIntegerRS_Qk_entry_0 ? 5'h0 : uIntergerRS_io_queue_data_split_0_qk; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_0_qk = uCDB_io_cdb_valid ? _GEN_2763 :
    uIntergerRS_io_queue_data_split_0_qk; 
  wire [131:0] uIntergerRS_io_update_entry_data_lo_lo = {uIntergerRS_io_queue_data_split_0_op,
    uIntergerRS_io_queue_data_split_0_dest,uIntergerRS_io_update_entry_data_split_0_qj,
    uIntergerRS_io_update_entry_data_split_0_qk,uIntergerRS_io_queue_data_split_0_a,
    uIntergerRS_io_update_entry_data_split_0_vj,uIntergerRS_io_update_entry_data_split_0_vk,
    uIntergerRS_io_queue_data_split_0_busy}; 
  wire [31:0] _GEN_2782 = need2_update_uIntegerRS_Qk_entry_1 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_1_vk
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_1_vk = uCDB_io_cdb_valid ? _GEN_2782 :
    uIntergerRS_io_queue_data_split_1_vk; 
  wire [31:0] _GEN_2780 = need2_update_uIntegerRS_Qj_entry_1 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_1_vj
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_1_vj = uCDB_io_cdb_valid ? _GEN_2780 :
    uIntergerRS_io_queue_data_split_1_vj; 
  wire [4:0] _GEN_2779 = need2_update_uIntegerRS_Qj_entry_1 ? 5'h0 : uIntergerRS_io_queue_data_split_1_qj; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_1_qj = uCDB_io_cdb_valid ? _GEN_2779 :
    uIntergerRS_io_queue_data_split_1_qj; 
  wire [4:0] _GEN_2781 = need2_update_uIntegerRS_Qk_entry_1 ? 5'h0 : uIntergerRS_io_queue_data_split_1_qk; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_1_qk = uCDB_io_cdb_valid ? _GEN_2781 :
    uIntergerRS_io_queue_data_split_1_qk; 
  wire [263:0] uIntergerRS_io_update_entry_data_lo = {uIntergerRS_io_queue_data_split_1_op,
    uIntergerRS_io_queue_data_split_1_dest,uIntergerRS_io_update_entry_data_split_1_qj,
    uIntergerRS_io_update_entry_data_split_1_qk,uIntergerRS_io_queue_data_split_1_a,
    uIntergerRS_io_update_entry_data_split_1_vj,uIntergerRS_io_update_entry_data_split_1_vk,
    uIntergerRS_io_queue_data_split_1_busy,uIntergerRS_io_update_entry_data_lo_lo}; 
  wire [31:0] _GEN_2800 = need2_update_uIntegerRS_Qk_entry_2 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_2_vk
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_2_vk = uCDB_io_cdb_valid ? _GEN_2800 :
    uIntergerRS_io_queue_data_split_2_vk; 
  wire [31:0] _GEN_2798 = need2_update_uIntegerRS_Qj_entry_2 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_2_vj
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_2_vj = uCDB_io_cdb_valid ? _GEN_2798 :
    uIntergerRS_io_queue_data_split_2_vj; 
  wire [4:0] _GEN_2797 = need2_update_uIntegerRS_Qj_entry_2 ? 5'h0 : uIntergerRS_io_queue_data_split_2_qj; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_2_qj = uCDB_io_cdb_valid ? _GEN_2797 :
    uIntergerRS_io_queue_data_split_2_qj; 
  wire [4:0] _GEN_2799 = need2_update_uIntegerRS_Qk_entry_2 ? 5'h0 : uIntergerRS_io_queue_data_split_2_qk; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_2_qk = uCDB_io_cdb_valid ? _GEN_2799 :
    uIntergerRS_io_queue_data_split_2_qk; 
  wire [131:0] uIntergerRS_io_update_entry_data_hi_lo = {uIntergerRS_io_queue_data_split_2_op,
    uIntergerRS_io_queue_data_split_2_dest,uIntergerRS_io_update_entry_data_split_2_qj,
    uIntergerRS_io_update_entry_data_split_2_qk,uIntergerRS_io_queue_data_split_2_a,
    uIntergerRS_io_update_entry_data_split_2_vj,uIntergerRS_io_update_entry_data_split_2_vk,
    uIntergerRS_io_queue_data_split_2_busy}; 
  wire [31:0] _GEN_2818 = need2_update_uIntegerRS_Qk_entry_3 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_3_vk
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_3_vk = uCDB_io_cdb_valid ? _GEN_2818 :
    uIntergerRS_io_queue_data_split_3_vk; 
  wire [31:0] _GEN_2816 = need2_update_uIntegerRS_Qj_entry_3 ? uCDB_io_cdb_result : uIntergerRS_io_queue_data_split_3_vj
    ; 
  wire [31:0] uIntergerRS_io_update_entry_data_split_3_vj = uCDB_io_cdb_valid ? _GEN_2816 :
    uIntergerRS_io_queue_data_split_3_vj; 
  wire [4:0] _GEN_2815 = need2_update_uIntegerRS_Qj_entry_3 ? 5'h0 : uIntergerRS_io_queue_data_split_3_qj; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_3_qj = uCDB_io_cdb_valid ? _GEN_2815 :
    uIntergerRS_io_queue_data_split_3_qj; 
  wire [4:0] _GEN_2817 = need2_update_uIntegerRS_Qk_entry_3 ? 5'h0 : uIntergerRS_io_queue_data_split_3_qk; 
  wire [4:0] uIntergerRS_io_update_entry_data_split_3_qk = uCDB_io_cdb_valid ? _GEN_2817 :
    uIntergerRS_io_queue_data_split_3_qk; 
  wire [263:0] uIntergerRS_io_update_entry_data_hi = {uIntergerRS_io_queue_data_split_3_op,
    uIntergerRS_io_queue_data_split_3_dest,uIntergerRS_io_update_entry_data_split_3_qj,
    uIntergerRS_io_update_entry_data_split_3_qk,uIntergerRS_io_queue_data_split_3_a,
    uIntergerRS_io_update_entry_data_split_3_vj,uIntergerRS_io_update_entry_data_split_3_vk,
    uIntergerRS_io_queue_data_split_3_busy,uIntergerRS_io_update_entry_data_hi_lo}; 
  wire  uMulDivRS_io_queue_data_split_0_busy = uMulDivRS__io_queue_data[0]; 
  wire [31:0] uMulDivRS_io_queue_data_split_0_vk = uMulDivRS__io_queue_data[32:1]; 
  wire [31:0] uMulDivRS_io_queue_data_split_0_vj = uMulDivRS__io_queue_data[64:33]; 
  wire [31:0] uMulDivRS_io_queue_data_split_0_a = uMulDivRS__io_queue_data[96:65]; 
  wire [4:0] uMulDivRS_io_queue_data_split_0_qk = uMulDivRS__io_queue_data[101:97]; 
  wire [4:0] uMulDivRS_io_queue_data_split_0_qj = uMulDivRS__io_queue_data[106:102]; 
  wire [4:0] uMulDivRS_io_queue_data_split_0_dest = uMulDivRS__io_queue_data[111:107]; 
  wire [19:0] uMulDivRS_io_queue_data_split_0_op = uMulDivRS__io_queue_data[131:112]; 
  wire  uMulDivRS_io_queue_data_split_1_busy = uMulDivRS__io_queue_data[132]; 
  wire [31:0] uMulDivRS_io_queue_data_split_1_vk = uMulDivRS__io_queue_data[164:133]; 
  wire [31:0] uMulDivRS_io_queue_data_split_1_vj = uMulDivRS__io_queue_data[196:165]; 
  wire [31:0] uMulDivRS_io_queue_data_split_1_a = uMulDivRS__io_queue_data[228:197]; 
  wire [4:0] uMulDivRS_io_queue_data_split_1_qk = uMulDivRS__io_queue_data[233:229]; 
  wire [4:0] uMulDivRS_io_queue_data_split_1_qj = uMulDivRS__io_queue_data[238:234]; 
  wire [4:0] uMulDivRS_io_queue_data_split_1_dest = uMulDivRS__io_queue_data[243:239]; 
  wire [19:0] uMulDivRS_io_queue_data_split_1_op = uMulDivRS__io_queue_data[263:244]; 
  wire  uMulDivRS_io_queue_data_split_2_busy = uMulDivRS__io_queue_data[264]; 
  wire [31:0] uMulDivRS_io_queue_data_split_2_vk = uMulDivRS__io_queue_data[296:265]; 
  wire [31:0] uMulDivRS_io_queue_data_split_2_vj = uMulDivRS__io_queue_data[328:297]; 
  wire [31:0] uMulDivRS_io_queue_data_split_2_a = uMulDivRS__io_queue_data[360:329]; 
  wire [4:0] uMulDivRS_io_queue_data_split_2_qk = uMulDivRS__io_queue_data[365:361]; 
  wire [4:0] uMulDivRS_io_queue_data_split_2_qj = uMulDivRS__io_queue_data[370:366]; 
  wire [4:0] uMulDivRS_io_queue_data_split_2_dest = uMulDivRS__io_queue_data[375:371]; 
  wire [19:0] uMulDivRS_io_queue_data_split_2_op = uMulDivRS__io_queue_data[395:376]; 
  wire  uMulDivRS_io_queue_data_split_3_busy = uMulDivRS__io_queue_data[396]; 
  wire [31:0] uMulDivRS_io_queue_data_split_3_vk = uMulDivRS__io_queue_data[428:397]; 
  wire [31:0] uMulDivRS_io_queue_data_split_3_vj = uMulDivRS__io_queue_data[460:429]; 
  wire [31:0] uMulDivRS_io_queue_data_split_3_a = uMulDivRS__io_queue_data[492:461]; 
  wire [4:0] uMulDivRS_io_queue_data_split_3_qk = uMulDivRS__io_queue_data[497:493]; 
  wire [4:0] uMulDivRS_io_queue_data_split_3_qj = uMulDivRS__io_queue_data[502:498]; 
  wire [4:0] uMulDivRS_io_queue_data_split_3_dest = uMulDivRS__io_queue_data[507:503]; 
  wire [19:0] uMulDivRS_io_queue_data_split_3_op = uMulDivRS__io_queue_data[527:508]; 
  wire [31:0] _GEN_2019 = ~uMulDivRS__io_full & _T_351 ? _GEN_422 : 32'h0; 
  wire [31:0] _GEN_2093 = muldiv_inst_r_io_d ? _GEN_2019 : 32'h0; 
  wire [31:0] _GEN_2240 = load_inst_r_io_d ? 32'h0 : _GEN_2093; 
  wire [31:0] _GEN_2323 = store_inst_r_io_d ? 32'h0 : _GEN_2240; 
  wire [31:0] _GEN_2413 = branch_inst_r_io_d ? 32'h0 : _GEN_2323; 
  wire [31:0] _GEN_2503 = integer_inst_r_io_d ? 32'h0 : _GEN_2413; 
  wire [31:0] uMulDivRS_io_enq_data_vk = decoder_if_inst_valid ? _GEN_2503 : 32'h0; 
  wire  _GEN_2085 = muldiv_inst_r_io_d & _T_409; 
  wire  _GEN_2235 = load_inst_r_io_d ? 1'h0 : _GEN_2085; 
  wire  _GEN_2318 = store_inst_r_io_d ? 1'h0 : _GEN_2235; 
  wire  _GEN_2408 = branch_inst_r_io_d ? 1'h0 : _GEN_2318; 
  wire  _GEN_2498 = integer_inst_r_io_d ? 1'h0 : _GEN_2408; 
  wire  uMulDivRS_io_enq_data_busy = decoder_if_inst_valid & _GEN_2498; 
  wire [31:0] _GEN_2017 = ~uMulDivRS__io_full & _T_351 ? _GEN_252 : 32'h0; 
  wire [31:0] _GEN_2091 = muldiv_inst_r_io_d ? _GEN_2017 : 32'h0; 
  wire [31:0] _GEN_2238 = load_inst_r_io_d ? 32'h0 : _GEN_2091; 
  wire [31:0] _GEN_2321 = store_inst_r_io_d ? 32'h0 : _GEN_2238; 
  wire [31:0] _GEN_2411 = branch_inst_r_io_d ? 32'h0 : _GEN_2321; 
  wire [31:0] _GEN_2501 = integer_inst_r_io_d ? 32'h0 : _GEN_2411; 
  wire [31:0] uMulDivRS_io_enq_data_vj = decoder_if_inst_valid ? _GEN_2501 : 32'h0; 
  wire [96:0] uMulDivRS_io_enq_data_lo = {32'h0,uMulDivRS_io_enq_data_vj,uMulDivRS_io_enq_data_vk,
    uMulDivRS_io_enq_data_busy}; 
  wire [4:0] _GEN_2018 = ~uMulDivRS__io_full & _T_351 ? _GEN_253 : 5'h0; 
  wire [4:0] _GEN_2092 = muldiv_inst_r_io_d ? _GEN_2018 : 5'h0; 
  wire [4:0] _GEN_2239 = load_inst_r_io_d ? 5'h0 : _GEN_2092; 
  wire [4:0] _GEN_2322 = store_inst_r_io_d ? 5'h0 : _GEN_2239; 
  wire [4:0] _GEN_2412 = branch_inst_r_io_d ? 5'h0 : _GEN_2322; 
  wire [4:0] _GEN_2502 = integer_inst_r_io_d ? 5'h0 : _GEN_2412; 
  wire [4:0] uMulDivRS_io_enq_data_qj = decoder_if_inst_valid ? _GEN_2502 : 5'h0; 
  wire [4:0] _GEN_2020 = ~uMulDivRS__io_full & _T_351 ? _GEN_423 : 5'h0; 
  wire [4:0] _GEN_2094 = muldiv_inst_r_io_d ? _GEN_2020 : 5'h0; 
  wire [4:0] _GEN_2241 = load_inst_r_io_d ? 5'h0 : _GEN_2094; 
  wire [4:0] _GEN_2324 = store_inst_r_io_d ? 5'h0 : _GEN_2241; 
  wire [4:0] _GEN_2414 = branch_inst_r_io_d ? 5'h0 : _GEN_2324; 
  wire [4:0] _GEN_2504 = integer_inst_r_io_d ? 5'h0 : _GEN_2414; 
  wire [4:0] uMulDivRS_io_enq_data_qk = decoder_if_inst_valid ? _GEN_2504 : 5'h0; 
  wire [19:0] _GEN_2015 = ~uMulDivRS__io_full & _T_351 ? _uIntergerRS_io_enq_data_op_T : 20'h0; 
  wire [19:0] _GEN_2089 = muldiv_inst_r_io_d ? _GEN_2015 : 20'h0; 
  wire [19:0] _GEN_2236 = load_inst_r_io_d ? 20'h0 : _GEN_2089; 
  wire [19:0] _GEN_2319 = store_inst_r_io_d ? 20'h0 : _GEN_2236; 
  wire [19:0] _GEN_2409 = branch_inst_r_io_d ? 20'h0 : _GEN_2319; 
  wire [19:0] _GEN_2499 = integer_inst_r_io_d ? 20'h0 : _GEN_2409; 
  wire [19:0] uMulDivRS_io_enq_data_op = decoder_if_inst_valid ? _GEN_2499 : 20'h0; 
  wire [4:0] _GEN_2016 = ~uMulDivRS__io_full & _T_351 ? uROB__io_enq_idx : 5'h0; 
  wire [4:0] _GEN_2090 = muldiv_inst_r_io_d ? _GEN_2016 : 5'h0; 
  wire [4:0] _GEN_2237 = load_inst_r_io_d ? 5'h0 : _GEN_2090; 
  wire [4:0] _GEN_2320 = store_inst_r_io_d ? 5'h0 : _GEN_2237; 
  wire [4:0] _GEN_2410 = branch_inst_r_io_d ? 5'h0 : _GEN_2320; 
  wire [4:0] _GEN_2500 = integer_inst_r_io_d ? 5'h0 : _GEN_2410; 
  wire [4:0] uMulDivRS_io_enq_data_dest = decoder_if_inst_valid ? _GEN_2500 : 5'h0; 
  wire [34:0] uMulDivRS_io_enq_data_hi = {uMulDivRS_io_enq_data_op,uMulDivRS_io_enq_data_dest,uMulDivRS_io_enq_data_qj,
    uMulDivRS_io_enq_data_qk}; 
  wire [4:0] uMulDivRS_io_deq_data_qk = uMulDivRS__io_deq_data[101:97]; 
  wire [4:0] uMulDivRS_io_deq_data_qj = uMulDivRS__io_deq_data[106:102]; 
  wire [19:0] uMulDivRS_io_deq_data_op = uMulDivRS__io_deq_data[131:112]; 
  wire  _T_566 = uMulDivRS_io_queue_data_split_1_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qj_entry_1 = _T_529 & _T_566; 
  wire  _T_568 = uMulDivRS_io_queue_data_split_1_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qk_entry_1 = _T_529 & _T_568; 
  wire  _T_570 = need2_update_uMulDivRS_Qj_entry_1 | need2_update_uMulDivRS_Qk_entry_1; 
  wire  uMulDivRS_io_update_entry_1 = _T_529 & _T_570; 
  wire  _T_557 = uMulDivRS_io_queue_data_split_0_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qj_entry_0 = _T_529 & _T_557; 
  wire  _T_559 = uMulDivRS_io_queue_data_split_0_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qk_entry_0 = _T_529 & _T_559; 
  wire  _T_561 = need2_update_uMulDivRS_Qj_entry_0 | need2_update_uMulDivRS_Qk_entry_0; 
  wire  uMulDivRS_io_update_entry_0 = _T_529 & _T_561; 
  wire [1:0] uMulDivRS_io_update_entry_lo = {uMulDivRS_io_update_entry_1,uMulDivRS_io_update_entry_0}; 
  wire  _T_584 = uMulDivRS_io_queue_data_split_3_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qj_entry_3 = _T_529 & _T_584; 
  wire  _T_586 = uMulDivRS_io_queue_data_split_3_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qk_entry_3 = _T_529 & _T_586; 
  wire  _T_588 = need2_update_uMulDivRS_Qj_entry_3 | need2_update_uMulDivRS_Qk_entry_3; 
  wire  uMulDivRS_io_update_entry_3 = _T_529 & _T_588; 
  wire  _T_575 = uMulDivRS_io_queue_data_split_2_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qj_entry_2 = _T_529 & _T_575; 
  wire  _T_577 = uMulDivRS_io_queue_data_split_2_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uMulDivRS_Qk_entry_2 = _T_529 & _T_577; 
  wire  _T_579 = need2_update_uMulDivRS_Qj_entry_2 | need2_update_uMulDivRS_Qk_entry_2; 
  wire  uMulDivRS_io_update_entry_2 = _T_529 & _T_579; 
  wire [1:0] uMulDivRS_io_update_entry_hi = {uMulDivRS_io_update_entry_3,uMulDivRS_io_update_entry_2}; 
  wire [31:0] _GEN_2836 = need2_update_uMulDivRS_Qk_entry_0 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_0_vk; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_0_vk = _T_529 ? _GEN_2836 : uMulDivRS_io_queue_data_split_0_vk; 
  wire [31:0] _GEN_2834 = need2_update_uMulDivRS_Qj_entry_0 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_0_vj; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_0_vj = _T_529 ? _GEN_2834 : uMulDivRS_io_queue_data_split_0_vj; 
  wire [4:0] _GEN_2833 = need2_update_uMulDivRS_Qj_entry_0 ? 5'h0 : uMulDivRS_io_queue_data_split_0_qj; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_0_qj = _T_529 ? _GEN_2833 : uMulDivRS_io_queue_data_split_0_qj; 
  wire [4:0] _GEN_2835 = need2_update_uMulDivRS_Qk_entry_0 ? 5'h0 : uMulDivRS_io_queue_data_split_0_qk; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_0_qk = _T_529 ? _GEN_2835 : uMulDivRS_io_queue_data_split_0_qk; 
  wire [131:0] uMulDivRS_io_update_entry_data_lo_lo = {uMulDivRS_io_queue_data_split_0_op,
    uMulDivRS_io_queue_data_split_0_dest,uMulDivRS_io_update_entry_data_split_0_qj,
    uMulDivRS_io_update_entry_data_split_0_qk,uMulDivRS_io_queue_data_split_0_a,
    uMulDivRS_io_update_entry_data_split_0_vj,uMulDivRS_io_update_entry_data_split_0_vk,
    uMulDivRS_io_queue_data_split_0_busy}; 
  wire [31:0] _GEN_2854 = need2_update_uMulDivRS_Qk_entry_1 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_1_vk; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_1_vk = _T_529 ? _GEN_2854 : uMulDivRS_io_queue_data_split_1_vk; 
  wire [31:0] _GEN_2852 = need2_update_uMulDivRS_Qj_entry_1 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_1_vj; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_1_vj = _T_529 ? _GEN_2852 : uMulDivRS_io_queue_data_split_1_vj; 
  wire [4:0] _GEN_2851 = need2_update_uMulDivRS_Qj_entry_1 ? 5'h0 : uMulDivRS_io_queue_data_split_1_qj; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_1_qj = _T_529 ? _GEN_2851 : uMulDivRS_io_queue_data_split_1_qj; 
  wire [4:0] _GEN_2853 = need2_update_uMulDivRS_Qk_entry_1 ? 5'h0 : uMulDivRS_io_queue_data_split_1_qk; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_1_qk = _T_529 ? _GEN_2853 : uMulDivRS_io_queue_data_split_1_qk; 
  wire [263:0] uMulDivRS_io_update_entry_data_lo = {uMulDivRS_io_queue_data_split_1_op,
    uMulDivRS_io_queue_data_split_1_dest,uMulDivRS_io_update_entry_data_split_1_qj,
    uMulDivRS_io_update_entry_data_split_1_qk,uMulDivRS_io_queue_data_split_1_a,
    uMulDivRS_io_update_entry_data_split_1_vj,uMulDivRS_io_update_entry_data_split_1_vk,
    uMulDivRS_io_queue_data_split_1_busy,uMulDivRS_io_update_entry_data_lo_lo}; 
  wire [31:0] _GEN_2872 = need2_update_uMulDivRS_Qk_entry_2 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_2_vk; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_2_vk = _T_529 ? _GEN_2872 : uMulDivRS_io_queue_data_split_2_vk; 
  wire [31:0] _GEN_2870 = need2_update_uMulDivRS_Qj_entry_2 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_2_vj; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_2_vj = _T_529 ? _GEN_2870 : uMulDivRS_io_queue_data_split_2_vj; 
  wire [4:0] _GEN_2869 = need2_update_uMulDivRS_Qj_entry_2 ? 5'h0 : uMulDivRS_io_queue_data_split_2_qj; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_2_qj = _T_529 ? _GEN_2869 : uMulDivRS_io_queue_data_split_2_qj; 
  wire [4:0] _GEN_2871 = need2_update_uMulDivRS_Qk_entry_2 ? 5'h0 : uMulDivRS_io_queue_data_split_2_qk; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_2_qk = _T_529 ? _GEN_2871 : uMulDivRS_io_queue_data_split_2_qk; 
  wire [131:0] uMulDivRS_io_update_entry_data_hi_lo = {uMulDivRS_io_queue_data_split_2_op,
    uMulDivRS_io_queue_data_split_2_dest,uMulDivRS_io_update_entry_data_split_2_qj,
    uMulDivRS_io_update_entry_data_split_2_qk,uMulDivRS_io_queue_data_split_2_a,
    uMulDivRS_io_update_entry_data_split_2_vj,uMulDivRS_io_update_entry_data_split_2_vk,
    uMulDivRS_io_queue_data_split_2_busy}; 
  wire [31:0] _GEN_2890 = need2_update_uMulDivRS_Qk_entry_3 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_3_vk; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_3_vk = _T_529 ? _GEN_2890 : uMulDivRS_io_queue_data_split_3_vk; 
  wire [31:0] _GEN_2888 = need2_update_uMulDivRS_Qj_entry_3 ? uCDB_io_cdb_result : uMulDivRS_io_queue_data_split_3_vj; 
  wire [31:0] uMulDivRS_io_update_entry_data_split_3_vj = _T_529 ? _GEN_2888 : uMulDivRS_io_queue_data_split_3_vj; 
  wire [4:0] _GEN_2887 = need2_update_uMulDivRS_Qj_entry_3 ? 5'h0 : uMulDivRS_io_queue_data_split_3_qj; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_3_qj = _T_529 ? _GEN_2887 : uMulDivRS_io_queue_data_split_3_qj; 
  wire [4:0] _GEN_2889 = need2_update_uMulDivRS_Qk_entry_3 ? 5'h0 : uMulDivRS_io_queue_data_split_3_qk; 
  wire [4:0] uMulDivRS_io_update_entry_data_split_3_qk = _T_529 ? _GEN_2889 : uMulDivRS_io_queue_data_split_3_qk; 
  wire [263:0] uMulDivRS_io_update_entry_data_hi = {uMulDivRS_io_queue_data_split_3_op,
    uMulDivRS_io_queue_data_split_3_dest,uMulDivRS_io_update_entry_data_split_3_qj,
    uMulDivRS_io_update_entry_data_split_3_qk,uMulDivRS_io_queue_data_split_3_a,
    uMulDivRS_io_update_entry_data_split_3_vj,uMulDivRS_io_update_entry_data_split_3_vk,
    uMulDivRS_io_queue_data_split_3_busy,uMulDivRS_io_update_entry_data_hi_lo}; 
  wire  uLoadStoreRS_io_queue_data_split_0_busy = uLoadStoreRS__io_queue_data[0]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_0_vk = uLoadStoreRS__io_queue_data[32:1]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_0_vj = uLoadStoreRS__io_queue_data[64:33]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_0_a = uLoadStoreRS__io_queue_data[96:65]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_0_qk = uLoadStoreRS__io_queue_data[101:97]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_0_qj = uLoadStoreRS__io_queue_data[106:102]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_0_dest = uLoadStoreRS__io_queue_data[111:107]; 
  wire [19:0] uLoadStoreRS_io_queue_data_split_0_op = uLoadStoreRS__io_queue_data[131:112]; 
  wire  uLoadStoreRS_io_queue_data_split_1_busy = uLoadStoreRS__io_queue_data[132]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_1_vk = uLoadStoreRS__io_queue_data[164:133]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_1_vj = uLoadStoreRS__io_queue_data[196:165]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_1_a = uLoadStoreRS__io_queue_data[228:197]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_1_qk = uLoadStoreRS__io_queue_data[233:229]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_1_qj = uLoadStoreRS__io_queue_data[238:234]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_1_dest = uLoadStoreRS__io_queue_data[243:239]; 
  wire [19:0] uLoadStoreRS_io_queue_data_split_1_op = uLoadStoreRS__io_queue_data[263:244]; 
  wire  uLoadStoreRS_io_queue_data_split_2_busy = uLoadStoreRS__io_queue_data[264]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_2_vk = uLoadStoreRS__io_queue_data[296:265]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_2_vj = uLoadStoreRS__io_queue_data[328:297]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_2_a = uLoadStoreRS__io_queue_data[360:329]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_2_qk = uLoadStoreRS__io_queue_data[365:361]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_2_qj = uLoadStoreRS__io_queue_data[370:366]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_2_dest = uLoadStoreRS__io_queue_data[375:371]; 
  wire [19:0] uLoadStoreRS_io_queue_data_split_2_op = uLoadStoreRS__io_queue_data[395:376]; 
  wire  uLoadStoreRS_io_queue_data_split_3_busy = uLoadStoreRS__io_queue_data[396]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_3_vk = uLoadStoreRS__io_queue_data[428:397]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_3_vj = uLoadStoreRS__io_queue_data[460:429]; 
  wire [31:0] uLoadStoreRS_io_queue_data_split_3_a = uLoadStoreRS__io_queue_data[492:461]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_3_qk = uLoadStoreRS__io_queue_data[497:493]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_3_qj = uLoadStoreRS__io_queue_data[502:498]; 
  wire [4:0] uLoadStoreRS_io_queue_data_split_3_dest = uLoadStoreRS__io_queue_data[507:503]; 
  wire [19:0] uLoadStoreRS_io_queue_data_split_3_op = uLoadStoreRS__io_queue_data[527:508]; 
  wire [31:0] _GEN_1264 = ~uLoadStoreRS__io_full & _T_351 ? _GEN_422 : 32'h0; 
  wire [31:0] _GEN_1541 = _T_384 ? _GEN_421 : 32'h0; 
  wire [31:0] _GEN_2169 = load_inst_r_io_d ? _GEN_1541 : 32'h0; 
  wire [31:0] _GEN_2252 = store_inst_r_io_d ? _GEN_1264 : _GEN_2169; 
  wire [31:0] _GEN_2342 = branch_inst_r_io_d ? 32'h0 : _GEN_2252; 
  wire [31:0] _GEN_2496 = integer_inst_r_io_d ? 32'h0 : _GEN_2342; 
  wire [31:0] uLoadStoreRS_io_enq_data_vk = decoder_if_inst_valid ? _GEN_2496 : 32'h0; 
  wire  _GEN_2163 = load_inst_r_io_d & _T_384; 
  wire  _GEN_2246 = store_inst_r_io_d ? _T_384 : _GEN_2163; 
  wire  _GEN_2336 = branch_inst_r_io_d ? 1'h0 : _GEN_2246; 
  wire  _GEN_2490 = integer_inst_r_io_d ? 1'h0 : _GEN_2336; 
  wire  uLoadStoreRS_io_enq_data_busy = decoder_if_inst_valid & _GEN_2490; 
  wire [31:0] _GEN_1261 = ~uLoadStoreRS__io_full & _T_351 ? decoder_if_imm : 32'h0; 
  wire [31:0] _GEN_2166 = load_inst_r_io_d ? _GEN_1261 : 32'h0; 
  wire [31:0] _GEN_2249 = store_inst_r_io_d ? _GEN_1261 : _GEN_2166; 
  wire [31:0] _GEN_2339 = branch_inst_r_io_d ? 32'h0 : _GEN_2249; 
  wire [31:0] _GEN_2493 = integer_inst_r_io_d ? 32'h0 : _GEN_2339; 
  wire [31:0] uLoadStoreRS_io_enq_data_a = decoder_if_inst_valid ? _GEN_2493 : 32'h0; 
  wire [31:0] _GEN_1262 = ~uLoadStoreRS__io_full & _T_351 ? _GEN_252 : 32'h0; 
  wire [31:0] _GEN_2167 = load_inst_r_io_d ? _GEN_1262 : 32'h0; 
  wire [31:0] _GEN_2250 = store_inst_r_io_d ? _GEN_1262 : _GEN_2167; 
  wire [31:0] _GEN_2340 = branch_inst_r_io_d ? 32'h0 : _GEN_2250; 
  wire [31:0] _GEN_2494 = integer_inst_r_io_d ? 32'h0 : _GEN_2340; 
  wire [31:0] uLoadStoreRS_io_enq_data_vj = decoder_if_inst_valid ? _GEN_2494 : 32'h0; 
  wire [96:0] uLoadStoreRS_io_enq_data_lo = {uLoadStoreRS_io_enq_data_a,uLoadStoreRS_io_enq_data_vj,
    uLoadStoreRS_io_enq_data_vk,uLoadStoreRS_io_enq_data_busy}; 
  wire [4:0] _GEN_1263 = ~uLoadStoreRS__io_full & _T_351 ? _GEN_253 : 5'h0; 
  wire [4:0] _GEN_2168 = load_inst_r_io_d ? _GEN_1263 : 5'h0; 
  wire [4:0] _GEN_2251 = store_inst_r_io_d ? _GEN_1263 : _GEN_2168; 
  wire [4:0] _GEN_2341 = branch_inst_r_io_d ? 5'h0 : _GEN_2251; 
  wire [4:0] _GEN_2495 = integer_inst_r_io_d ? 5'h0 : _GEN_2341; 
  wire [4:0] uLoadStoreRS_io_enq_data_qj = decoder_if_inst_valid ? _GEN_2495 : 5'h0; 
  wire [4:0] _GEN_1265 = ~uLoadStoreRS__io_full & _T_351 ? _GEN_423 : 5'h0; 
  wire [4:0] _GEN_2253 = store_inst_r_io_d ? _GEN_1265 : 5'h0; 
  wire [4:0] _GEN_2343 = branch_inst_r_io_d ? 5'h0 : _GEN_2253; 
  wire [4:0] _GEN_2497 = integer_inst_r_io_d ? 5'h0 : _GEN_2343; 
  wire [4:0] uLoadStoreRS_io_enq_data_qk = decoder_if_inst_valid ? _GEN_2497 : 5'h0; 
  wire [19:0] _GEN_1259 = ~uLoadStoreRS__io_full & _T_351 ? _uIntergerRS_io_enq_data_op_T : 20'h0; 
  wire [19:0] _GEN_2164 = load_inst_r_io_d ? _GEN_1259 : 20'h0; 
  wire [19:0] _GEN_2247 = store_inst_r_io_d ? _GEN_1259 : _GEN_2164; 
  wire [19:0] _GEN_2337 = branch_inst_r_io_d ? 20'h0 : _GEN_2247; 
  wire [19:0] _GEN_2491 = integer_inst_r_io_d ? 20'h0 : _GEN_2337; 
  wire [19:0] uLoadStoreRS_io_enq_data_op = decoder_if_inst_valid ? _GEN_2491 : 20'h0; 
  wire [4:0] _GEN_1260 = ~uLoadStoreRS__io_full & _T_351 ? uROB__io_enq_idx : 5'h0; 
  wire [4:0] _GEN_2165 = load_inst_r_io_d ? _GEN_1260 : 5'h0; 
  wire [4:0] _GEN_2248 = store_inst_r_io_d ? _GEN_1260 : _GEN_2165; 
  wire [4:0] _GEN_2338 = branch_inst_r_io_d ? 5'h0 : _GEN_2248; 
  wire [4:0] _GEN_2492 = integer_inst_r_io_d ? 5'h0 : _GEN_2338; 
  wire [4:0] uLoadStoreRS_io_enq_data_dest = decoder_if_inst_valid ? _GEN_2492 : 5'h0; 
  wire [34:0] uLoadStoreRS_io_enq_data_hi = {uLoadStoreRS_io_enq_data_op,uLoadStoreRS_io_enq_data_dest,
    uLoadStoreRS_io_enq_data_qj,uLoadStoreRS_io_enq_data_qk}; 
  wire  _T_602 = uLoadStoreRS_io_queue_data_split_1_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qj_entry_1 = _T_529 & _T_602; 
  wire  _T_604 = uLoadStoreRS_io_queue_data_split_1_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qk_entry_1 = _T_529 & _T_604; 
  wire  _T_606 = need2_update_uLoadStoreRS_Qj_entry_1 | need2_update_uLoadStoreRS_Qk_entry_1; 
  wire  uLoadStoreRS_io_update_entry_1 = _T_529 & _T_606; 
  wire  _T_593 = uLoadStoreRS_io_queue_data_split_0_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qj_entry_0 = _T_529 & _T_593; 
  wire  _T_595 = uLoadStoreRS_io_queue_data_split_0_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qk_entry_0 = _T_529 & _T_595; 
  wire  _T_597 = need2_update_uLoadStoreRS_Qj_entry_0 | need2_update_uLoadStoreRS_Qk_entry_0; 
  wire  uLoadStoreRS_io_update_entry_0 = _T_529 & _T_597; 
  wire [1:0] uLoadStoreRS_io_update_entry_lo = {uLoadStoreRS_io_update_entry_1,uLoadStoreRS_io_update_entry_0}; 
  wire  _T_620 = uLoadStoreRS_io_queue_data_split_3_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qj_entry_3 = _T_529 & _T_620; 
  wire  _T_622 = uLoadStoreRS_io_queue_data_split_3_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qk_entry_3 = _T_529 & _T_622; 
  wire  _T_624 = need2_update_uLoadStoreRS_Qj_entry_3 | need2_update_uLoadStoreRS_Qk_entry_3; 
  wire  uLoadStoreRS_io_update_entry_3 = _T_529 & _T_624; 
  wire  _T_611 = uLoadStoreRS_io_queue_data_split_2_qj == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qj_entry_2 = _T_529 & _T_611; 
  wire  _T_613 = uLoadStoreRS_io_queue_data_split_2_qk == uCDB_io_cdb_dest; 
  wire  need2_update_uLoadStoreRS_Qk_entry_2 = _T_529 & _T_613; 
  wire  _T_615 = need2_update_uLoadStoreRS_Qj_entry_2 | need2_update_uLoadStoreRS_Qk_entry_2; 
  wire  uLoadStoreRS_io_update_entry_2 = _T_529 & _T_615; 
  wire [1:0] uLoadStoreRS_io_update_entry_hi = {uLoadStoreRS_io_update_entry_3,uLoadStoreRS_io_update_entry_2}; 
  wire [31:0] _GEN_2908 = need2_update_uLoadStoreRS_Qk_entry_0 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_0_vk; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_0_vk = _T_529 ? _GEN_2908 : uLoadStoreRS_io_queue_data_split_0_vk; 
  wire [31:0] _GEN_2906 = need2_update_uLoadStoreRS_Qj_entry_0 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_0_vj; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_0_vj = _T_529 ? _GEN_2906 : uLoadStoreRS_io_queue_data_split_0_vj; 
  wire [4:0] _GEN_2905 = need2_update_uLoadStoreRS_Qj_entry_0 ? 5'h0 : uLoadStoreRS_io_queue_data_split_0_qj; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_0_qj = _T_529 ? _GEN_2905 : uLoadStoreRS_io_queue_data_split_0_qj; 
  wire [4:0] _GEN_2907 = need2_update_uLoadStoreRS_Qk_entry_0 ? 5'h0 : uLoadStoreRS_io_queue_data_split_0_qk; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_0_qk = _T_529 ? _GEN_2907 : uLoadStoreRS_io_queue_data_split_0_qk; 
  wire [131:0] uLoadStoreRS_io_update_entry_data_lo_lo = {uLoadStoreRS_io_queue_data_split_0_op,
    uLoadStoreRS_io_queue_data_split_0_dest,uLoadStoreRS_io_update_entry_data_split_0_qj,
    uLoadStoreRS_io_update_entry_data_split_0_qk,uLoadStoreRS_io_queue_data_split_0_a,
    uLoadStoreRS_io_update_entry_data_split_0_vj,uLoadStoreRS_io_update_entry_data_split_0_vk,
    uLoadStoreRS_io_queue_data_split_0_busy}; 
  wire [31:0] _GEN_2926 = need2_update_uLoadStoreRS_Qk_entry_1 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_1_vk; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_1_vk = _T_529 ? _GEN_2926 : uLoadStoreRS_io_queue_data_split_1_vk; 
  wire [31:0] _GEN_2924 = need2_update_uLoadStoreRS_Qj_entry_1 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_1_vj; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_1_vj = _T_529 ? _GEN_2924 : uLoadStoreRS_io_queue_data_split_1_vj; 
  wire [4:0] _GEN_2923 = need2_update_uLoadStoreRS_Qj_entry_1 ? 5'h0 : uLoadStoreRS_io_queue_data_split_1_qj; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_1_qj = _T_529 ? _GEN_2923 : uLoadStoreRS_io_queue_data_split_1_qj; 
  wire [4:0] _GEN_2925 = need2_update_uLoadStoreRS_Qk_entry_1 ? 5'h0 : uLoadStoreRS_io_queue_data_split_1_qk; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_1_qk = _T_529 ? _GEN_2925 : uLoadStoreRS_io_queue_data_split_1_qk; 
  wire [263:0] uLoadStoreRS_io_update_entry_data_lo = {uLoadStoreRS_io_queue_data_split_1_op,
    uLoadStoreRS_io_queue_data_split_1_dest,uLoadStoreRS_io_update_entry_data_split_1_qj,
    uLoadStoreRS_io_update_entry_data_split_1_qk,uLoadStoreRS_io_queue_data_split_1_a,
    uLoadStoreRS_io_update_entry_data_split_1_vj,uLoadStoreRS_io_update_entry_data_split_1_vk,
    uLoadStoreRS_io_queue_data_split_1_busy,uLoadStoreRS_io_update_entry_data_lo_lo}; 
  wire [31:0] _GEN_2944 = need2_update_uLoadStoreRS_Qk_entry_2 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_2_vk; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_2_vk = _T_529 ? _GEN_2944 : uLoadStoreRS_io_queue_data_split_2_vk; 
  wire [31:0] _GEN_2942 = need2_update_uLoadStoreRS_Qj_entry_2 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_2_vj; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_2_vj = _T_529 ? _GEN_2942 : uLoadStoreRS_io_queue_data_split_2_vj; 
  wire [4:0] _GEN_2941 = need2_update_uLoadStoreRS_Qj_entry_2 ? 5'h0 : uLoadStoreRS_io_queue_data_split_2_qj; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_2_qj = _T_529 ? _GEN_2941 : uLoadStoreRS_io_queue_data_split_2_qj; 
  wire [4:0] _GEN_2943 = need2_update_uLoadStoreRS_Qk_entry_2 ? 5'h0 : uLoadStoreRS_io_queue_data_split_2_qk; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_2_qk = _T_529 ? _GEN_2943 : uLoadStoreRS_io_queue_data_split_2_qk; 
  wire [131:0] uLoadStoreRS_io_update_entry_data_hi_lo = {uLoadStoreRS_io_queue_data_split_2_op,
    uLoadStoreRS_io_queue_data_split_2_dest,uLoadStoreRS_io_update_entry_data_split_2_qj,
    uLoadStoreRS_io_update_entry_data_split_2_qk,uLoadStoreRS_io_queue_data_split_2_a,
    uLoadStoreRS_io_update_entry_data_split_2_vj,uLoadStoreRS_io_update_entry_data_split_2_vk,
    uLoadStoreRS_io_queue_data_split_2_busy}; 
  wire [31:0] _GEN_2962 = need2_update_uLoadStoreRS_Qk_entry_3 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_3_vk; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_3_vk = _T_529 ? _GEN_2962 : uLoadStoreRS_io_queue_data_split_3_vk; 
  wire [31:0] _GEN_2960 = need2_update_uLoadStoreRS_Qj_entry_3 ? uCDB_io_cdb_result :
    uLoadStoreRS_io_queue_data_split_3_vj; 
  wire [31:0] uLoadStoreRS_io_update_entry_data_split_3_vj = _T_529 ? _GEN_2960 : uLoadStoreRS_io_queue_data_split_3_vj; 
  wire [4:0] _GEN_2959 = need2_update_uLoadStoreRS_Qj_entry_3 ? 5'h0 : uLoadStoreRS_io_queue_data_split_3_qj; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_3_qj = _T_529 ? _GEN_2959 : uLoadStoreRS_io_queue_data_split_3_qj; 
  wire [4:0] _GEN_2961 = need2_update_uLoadStoreRS_Qk_entry_3 ? 5'h0 : uLoadStoreRS_io_queue_data_split_3_qk; 
  wire [4:0] uLoadStoreRS_io_update_entry_data_split_3_qk = _T_529 ? _GEN_2961 : uLoadStoreRS_io_queue_data_split_3_qk; 
  wire [263:0] uLoadStoreRS_io_update_entry_data_hi = {uLoadStoreRS_io_queue_data_split_3_op,
    uLoadStoreRS_io_queue_data_split_3_dest,uLoadStoreRS_io_update_entry_data_split_3_qj,
    uLoadStoreRS_io_update_entry_data_split_3_qk,uLoadStoreRS_io_queue_data_split_3_a,
    uLoadStoreRS_io_update_entry_data_split_3_vj,uLoadStoreRS_io_update_entry_data_split_3_vk,
    uLoadStoreRS_io_queue_data_split_3_busy,uLoadStoreRS_io_update_entry_data_hi_lo}; 
  wire [1:0] branchProc_stEnum = mBranchProc_st_io_q; 
  wire  _integer_inst_r_io_d_T = decoder_if_exe_op_and | decoder_if_exe_op_or; 
  wire  _integer_inst_r_io_d_T_1 = _integer_inst_r_io_d_T | decoder_if_exe_op_xor; 
  wire  _integer_inst_r_io_d_T_2 = _integer_inst_r_io_d_T_1 | decoder_if_exe_op_set; 
  wire  _integer_inst_r_io_d_T_3 = _integer_inst_r_io_d_T_2 | decoder_if_exe_op_add; 
  wire  _integer_inst_r_io_d_T_4 = _integer_inst_r_io_d_T_3 | decoder_if_exe_op_sub; 
  wire  _integer_inst_r_io_d_T_5 = _integer_inst_r_io_d_T_4 | decoder_if_exe_op_sll; 
  wire  _integer_inst_r_io_d_T_6 = _integer_inst_r_io_d_T_5 | decoder_if_exe_op_srl; 
  wire  _integer_inst_r_io_d_T_7 = _integer_inst_r_io_d_T_6 | decoder_if_exe_op_sra; 
  wire  _integer_inst_r_io_d_T_8 = ~decoder_if_exe_op_br; 
  wire  _integer_inst_r_io_d_T_9 = ~decoder_if_exe_op_br & decoder_if_exe_op_less; 
  wire  _integer_inst_r_io_d_T_10 = _integer_inst_r_io_d_T_7 | _integer_inst_r_io_d_T_9; 
  wire  _integer_inst_r_io_d_T_12 = _integer_inst_r_io_d_T_8 & decoder_if_exe_op_large; 
  wire  _integer_inst_r_io_d_T_13 = _integer_inst_r_io_d_T_10 | _integer_inst_r_io_d_T_12; 
  wire  _integer_inst_r_io_d_T_15 = _integer_inst_r_io_d_T_8 & decoder_if_exe_op_equal; 
  wire  _T_39 = uIntergerRS__io_full | uROB__io_full; 
  wire [1:0] _GEN_1 = uIntergerRS__io_full | uROB__io_full ? 2'h1 : mBranchProc_st_io_q; 
  wire  _T_43 = uLoadStoreRS__io_full | uROB__io_full; 
  wire [1:0] _GEN_3 = uLoadStoreRS__io_full | uROB__io_full ? 2'h1 : mBranchProc_st_io_q; 
  wire  _T_46 = uMulDivRS__io_full | uROB__io_full; 
  wire [1:0] _GEN_5 = uMulDivRS__io_full | uROB__io_full ? 2'h1 : mBranchProc_st_io_q; 
  wire  _GEN_6 = _T_406 & _T_46; 
  wire [1:0] _GEN_7 = _T_406 ? _GEN_5 : mBranchProc_st_io_q; 
  wire  _GEN_8 = store_inst_r_io_d | load_inst_r_io_d ? _T_43 : _GEN_6; 
  wire [1:0] _GEN_9 = store_inst_r_io_d | load_inst_r_io_d ? _GEN_3 : _GEN_7; 
  wire  _GEN_10 = integer_inst_r_io_d | branch_inst_r_io_d ? _T_39 : _GEN_8; 
  wire [1:0] _GEN_11 = integer_inst_r_io_d | branch_inst_r_io_d ? _GEN_1 : _GEN_9; 
  wire  _GEN_12 = decoder_if_inst_valid & _GEN_10; 
  wire [1:0] _GEN_13 = decoder_if_inst_valid ? _GEN_11 : mBranchProc_st_io_q; 
  wire  _T_52 = uIntergerRS__io_full & (integer_inst_r_io_q | branch_inst_r_io_q); 
  wire  _T_53 = uROB__io_full | _T_52; 
  wire  _T_55 = uLoadStoreRS__io_full & (store_inst_r_io_q | load_inst_r_io_q); 
  wire  _T_56 = _T_53 | _T_55; 
  wire  _T_57 = uMulDivRS__io_full & muldiv_inst_r_io_q; 
  wire  _T_58 = _T_56 | _T_57; 
  wire  _GEN_16 = 2'h1 == branchProc_stEnum & _T_58; 
  wire [1:0] _GEN_17 = 2'h1 == branchProc_stEnum ? {{1'd0}, _T_58} : mBranchProc_st_io_q; 
  wire  _T_61 = uROB_io_deq_data_rob_type == 2'h1; 
  wire  _T_62 = uROB__io_deq & _T_61; 
  wire  _T_64 = 5'h0 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_65 = _T_62 & _T_64; 
  wire  _T_66 = uRegState_io_0_q_reorder == uROB__io_deq_idx; 
  wire  _T_67 = _T_65 & _T_66; 
  wire [4:0] _GEN_20 = _T_67 ? 5'h0 : uRegState_io_0_q_reorder; 
  wire  _GEN_21 = _T_67 ? 1'h0 : uRegState_io_0_q_busy; 
  wire  _T_73 = 5'h1 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_74 = _T_62 & _T_73; 
  wire  _T_75 = uRegState_io_1_q_reorder == uROB__io_deq_idx; 
  wire  _T_76 = _T_74 & _T_75; 
  wire [4:0] _GEN_22 = _T_76 ? 5'h0 : uRegState_io_1_q_reorder; 
  wire  _GEN_23 = _T_76 ? 1'h0 : uRegState_io_1_q_busy; 
  wire  _T_82 = 5'h2 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_83 = _T_62 & _T_82; 
  wire  _T_84 = uRegState_io_2_q_reorder == uROB__io_deq_idx; 
  wire  _T_85 = _T_83 & _T_84; 
  wire [4:0] _GEN_24 = _T_85 ? 5'h0 : uRegState_io_2_q_reorder; 
  wire  _GEN_25 = _T_85 ? 1'h0 : uRegState_io_2_q_busy; 
  wire  _T_91 = 5'h3 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_92 = _T_62 & _T_91; 
  wire  _T_93 = uRegState_io_3_q_reorder == uROB__io_deq_idx; 
  wire  _T_94 = _T_92 & _T_93; 
  wire [4:0] _GEN_26 = _T_94 ? 5'h0 : uRegState_io_3_q_reorder; 
  wire  _GEN_27 = _T_94 ? 1'h0 : uRegState_io_3_q_busy; 
  wire  _T_100 = 5'h4 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_101 = _T_62 & _T_100; 
  wire  _T_102 = uRegState_io_4_q_reorder == uROB__io_deq_idx; 
  wire  _T_103 = _T_101 & _T_102; 
  wire [4:0] _GEN_28 = _T_103 ? 5'h0 : uRegState_io_4_q_reorder; 
  wire  _GEN_29 = _T_103 ? 1'h0 : uRegState_io_4_q_busy; 
  wire  _T_109 = 5'h5 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_110 = _T_62 & _T_109; 
  wire  _T_111 = uRegState_io_5_q_reorder == uROB__io_deq_idx; 
  wire  _T_112 = _T_110 & _T_111; 
  wire [4:0] _GEN_30 = _T_112 ? 5'h0 : uRegState_io_5_q_reorder; 
  wire  _GEN_31 = _T_112 ? 1'h0 : uRegState_io_5_q_busy; 
  wire  _T_118 = 5'h6 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_119 = _T_62 & _T_118; 
  wire  _T_120 = uRegState_io_6_q_reorder == uROB__io_deq_idx; 
  wire  _T_121 = _T_119 & _T_120; 
  wire [4:0] _GEN_32 = _T_121 ? 5'h0 : uRegState_io_6_q_reorder; 
  wire  _GEN_33 = _T_121 ? 1'h0 : uRegState_io_6_q_busy; 
  wire  _T_127 = 5'h7 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_128 = _T_62 & _T_127; 
  wire  _T_129 = uRegState_io_7_q_reorder == uROB__io_deq_idx; 
  wire  _T_130 = _T_128 & _T_129; 
  wire [4:0] _GEN_34 = _T_130 ? 5'h0 : uRegState_io_7_q_reorder; 
  wire  _GEN_35 = _T_130 ? 1'h0 : uRegState_io_7_q_busy; 
  wire  _T_136 = 5'h8 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_137 = _T_62 & _T_136; 
  wire  _T_138 = uRegState_io_8_q_reorder == uROB__io_deq_idx; 
  wire  _T_139 = _T_137 & _T_138; 
  wire [4:0] _GEN_36 = _T_139 ? 5'h0 : uRegState_io_8_q_reorder; 
  wire  _GEN_37 = _T_139 ? 1'h0 : uRegState_io_8_q_busy; 
  wire  _T_145 = 5'h9 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_146 = _T_62 & _T_145; 
  wire  _T_147 = uRegState_io_9_q_reorder == uROB__io_deq_idx; 
  wire  _T_148 = _T_146 & _T_147; 
  wire [4:0] _GEN_38 = _T_148 ? 5'h0 : uRegState_io_9_q_reorder; 
  wire  _GEN_39 = _T_148 ? 1'h0 : uRegState_io_9_q_busy; 
  wire  _T_154 = 5'ha == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_155 = _T_62 & _T_154; 
  wire  _T_156 = uRegState_io_10_q_reorder == uROB__io_deq_idx; 
  wire  _T_157 = _T_155 & _T_156; 
  wire [4:0] _GEN_40 = _T_157 ? 5'h0 : uRegState_io_10_q_reorder; 
  wire  _GEN_41 = _T_157 ? 1'h0 : uRegState_io_10_q_busy; 
  wire  _T_163 = 5'hb == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_164 = _T_62 & _T_163; 
  wire  _T_165 = uRegState_io_11_q_reorder == uROB__io_deq_idx; 
  wire  _T_166 = _T_164 & _T_165; 
  wire [4:0] _GEN_42 = _T_166 ? 5'h0 : uRegState_io_11_q_reorder; 
  wire  _GEN_43 = _T_166 ? 1'h0 : uRegState_io_11_q_busy; 
  wire  _T_172 = 5'hc == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_173 = _T_62 & _T_172; 
  wire  _T_174 = uRegState_io_12_q_reorder == uROB__io_deq_idx; 
  wire  _T_175 = _T_173 & _T_174; 
  wire [4:0] _GEN_44 = _T_175 ? 5'h0 : uRegState_io_12_q_reorder; 
  wire  _GEN_45 = _T_175 ? 1'h0 : uRegState_io_12_q_busy; 
  wire  _T_181 = 5'hd == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_182 = _T_62 & _T_181; 
  wire  _T_183 = uRegState_io_13_q_reorder == uROB__io_deq_idx; 
  wire  _T_184 = _T_182 & _T_183; 
  wire [4:0] _GEN_46 = _T_184 ? 5'h0 : uRegState_io_13_q_reorder; 
  wire  _GEN_47 = _T_184 ? 1'h0 : uRegState_io_13_q_busy; 
  wire  _T_190 = 5'he == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_191 = _T_62 & _T_190; 
  wire  _T_192 = uRegState_io_14_q_reorder == uROB__io_deq_idx; 
  wire  _T_193 = _T_191 & _T_192; 
  wire [4:0] _GEN_48 = _T_193 ? 5'h0 : uRegState_io_14_q_reorder; 
  wire  _GEN_49 = _T_193 ? 1'h0 : uRegState_io_14_q_busy; 
  wire  _T_199 = 5'hf == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_200 = _T_62 & _T_199; 
  wire  _T_201 = uRegState_io_15_q_reorder == uROB__io_deq_idx; 
  wire  _T_202 = _T_200 & _T_201; 
  wire [4:0] _GEN_50 = _T_202 ? 5'h0 : uRegState_io_15_q_reorder; 
  wire  _GEN_51 = _T_202 ? 1'h0 : uRegState_io_15_q_busy; 
  wire  _T_208 = 5'h10 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_209 = _T_62 & _T_208; 
  wire  _T_210 = uRegState_io_16_q_reorder == uROB__io_deq_idx; 
  wire  _T_211 = _T_209 & _T_210; 
  wire [4:0] _GEN_52 = _T_211 ? 5'h0 : uRegState_io_16_q_reorder; 
  wire  _GEN_53 = _T_211 ? 1'h0 : uRegState_io_16_q_busy; 
  wire  _T_217 = 5'h11 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_218 = _T_62 & _T_217; 
  wire  _T_219 = uRegState_io_17_q_reorder == uROB__io_deq_idx; 
  wire  _T_220 = _T_218 & _T_219; 
  wire [4:0] _GEN_54 = _T_220 ? 5'h0 : uRegState_io_17_q_reorder; 
  wire  _GEN_55 = _T_220 ? 1'h0 : uRegState_io_17_q_busy; 
  wire  _T_226 = 5'h12 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_227 = _T_62 & _T_226; 
  wire  _T_228 = uRegState_io_18_q_reorder == uROB__io_deq_idx; 
  wire  _T_229 = _T_227 & _T_228; 
  wire [4:0] _GEN_56 = _T_229 ? 5'h0 : uRegState_io_18_q_reorder; 
  wire  _GEN_57 = _T_229 ? 1'h0 : uRegState_io_18_q_busy; 
  wire  _T_235 = 5'h13 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_236 = _T_62 & _T_235; 
  wire  _T_237 = uRegState_io_19_q_reorder == uROB__io_deq_idx; 
  wire  _T_238 = _T_236 & _T_237; 
  wire [4:0] _GEN_58 = _T_238 ? 5'h0 : uRegState_io_19_q_reorder; 
  wire  _GEN_59 = _T_238 ? 1'h0 : uRegState_io_19_q_busy; 
  wire  _T_244 = 5'h14 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_245 = _T_62 & _T_244; 
  wire  _T_246 = uRegState_io_20_q_reorder == uROB__io_deq_idx; 
  wire  _T_247 = _T_245 & _T_246; 
  wire [4:0] _GEN_60 = _T_247 ? 5'h0 : uRegState_io_20_q_reorder; 
  wire  _GEN_61 = _T_247 ? 1'h0 : uRegState_io_20_q_busy; 
  wire  _T_253 = 5'h15 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_254 = _T_62 & _T_253; 
  wire  _T_255 = uRegState_io_21_q_reorder == uROB__io_deq_idx; 
  wire  _T_256 = _T_254 & _T_255; 
  wire [4:0] _GEN_62 = _T_256 ? 5'h0 : uRegState_io_21_q_reorder; 
  wire  _GEN_63 = _T_256 ? 1'h0 : uRegState_io_21_q_busy; 
  wire  _T_262 = 5'h16 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_263 = _T_62 & _T_262; 
  wire  _T_264 = uRegState_io_22_q_reorder == uROB__io_deq_idx; 
  wire  _T_265 = _T_263 & _T_264; 
  wire [4:0] _GEN_64 = _T_265 ? 5'h0 : uRegState_io_22_q_reorder; 
  wire  _GEN_65 = _T_265 ? 1'h0 : uRegState_io_22_q_busy; 
  wire  _T_271 = 5'h17 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_272 = _T_62 & _T_271; 
  wire  _T_273 = uRegState_io_23_q_reorder == uROB__io_deq_idx; 
  wire  _T_274 = _T_272 & _T_273; 
  wire [4:0] _GEN_66 = _T_274 ? 5'h0 : uRegState_io_23_q_reorder; 
  wire  _GEN_67 = _T_274 ? 1'h0 : uRegState_io_23_q_busy; 
  wire  _T_280 = 5'h18 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_281 = _T_62 & _T_280; 
  wire  _T_282 = uRegState_io_24_q_reorder == uROB__io_deq_idx; 
  wire  _T_283 = _T_281 & _T_282; 
  wire [4:0] _GEN_68 = _T_283 ? 5'h0 : uRegState_io_24_q_reorder; 
  wire  _GEN_69 = _T_283 ? 1'h0 : uRegState_io_24_q_busy; 
  wire  _T_289 = 5'h19 == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_290 = _T_62 & _T_289; 
  wire  _T_291 = uRegState_io_25_q_reorder == uROB__io_deq_idx; 
  wire  _T_292 = _T_290 & _T_291; 
  wire [4:0] _GEN_70 = _T_292 ? 5'h0 : uRegState_io_25_q_reorder; 
  wire  _GEN_71 = _T_292 ? 1'h0 : uRegState_io_25_q_busy; 
  wire  _T_298 = 5'h1a == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_299 = _T_62 & _T_298; 
  wire  _T_300 = uRegState_io_26_q_reorder == uROB__io_deq_idx; 
  wire  _T_301 = _T_299 & _T_300; 
  wire [4:0] _GEN_72 = _T_301 ? 5'h0 : uRegState_io_26_q_reorder; 
  wire  _GEN_73 = _T_301 ? 1'h0 : uRegState_io_26_q_busy; 
  wire  _T_307 = 5'h1b == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_308 = _T_62 & _T_307; 
  wire  _T_309 = uRegState_io_27_q_reorder == uROB__io_deq_idx; 
  wire  _T_310 = _T_308 & _T_309; 
  wire [4:0] _GEN_74 = _T_310 ? 5'h0 : uRegState_io_27_q_reorder; 
  wire  _GEN_75 = _T_310 ? 1'h0 : uRegState_io_27_q_busy; 
  wire  _T_316 = 5'h1c == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_317 = _T_62 & _T_316; 
  wire  _T_318 = uRegState_io_28_q_reorder == uROB__io_deq_idx; 
  wire  _T_319 = _T_317 & _T_318; 
  wire [4:0] _GEN_76 = _T_319 ? 5'h0 : uRegState_io_28_q_reorder; 
  wire  _GEN_77 = _T_319 ? 1'h0 : uRegState_io_28_q_busy; 
  wire  _T_325 = 5'h1d == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_326 = _T_62 & _T_325; 
  wire  _T_327 = uRegState_io_29_q_reorder == uROB__io_deq_idx; 
  wire  _T_328 = _T_326 & _T_327; 
  wire [4:0] _GEN_78 = _T_328 ? 5'h0 : uRegState_io_29_q_reorder; 
  wire  _GEN_79 = _T_328 ? 1'h0 : uRegState_io_29_q_busy; 
  wire  _T_334 = 5'h1e == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_335 = _T_62 & _T_334; 
  wire  _T_336 = uRegState_io_30_q_reorder == uROB__io_deq_idx; 
  wire  _T_337 = _T_335 & _T_336; 
  wire [4:0] _GEN_80 = _T_337 ? 5'h0 : uRegState_io_30_q_reorder; 
  wire  _GEN_81 = _T_337 ? 1'h0 : uRegState_io_30_q_busy; 
  wire  _T_343 = 5'h1f == uROB_io_deq_data_rob_dest[4:0]; 
  wire  _T_344 = _T_62 & _T_343; 
  wire  _T_345 = uRegState_io_31_q_reorder == uROB__io_deq_idx; 
  wire  _T_346 = _T_344 & _T_345; 
  wire [4:0] _GEN_82 = _T_346 ? 5'h0 : uRegState_io_31_q_reorder; 
  wire  _GEN_83 = _T_346 ? 1'h0 : uRegState_io_31_q_busy; 
  wire [4:0] _uRegState_io_decoder_if_rd_idx_d_reorder = uROB__io_enq_idx; 
  wire [4:0] _GEN_427 = 5'h0 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_20; 
  wire [4:0] _GEN_428 = 5'h1 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_22; 
  wire [4:0] _GEN_429 = 5'h2 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_24; 
  wire [4:0] _GEN_430 = 5'h3 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_26; 
  wire [4:0] _GEN_431 = 5'h4 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_28; 
  wire [4:0] _GEN_432 = 5'h5 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_30; 
  wire [4:0] _GEN_433 = 5'h6 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_32; 
  wire [4:0] _GEN_434 = 5'h7 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_34; 
  wire [4:0] _GEN_435 = 5'h8 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_36; 
  wire [4:0] _GEN_436 = 5'h9 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_38; 
  wire [4:0] _GEN_437 = 5'ha == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_40; 
  wire [4:0] _GEN_438 = 5'hb == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_42; 
  wire [4:0] _GEN_439 = 5'hc == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_44; 
  wire [4:0] _GEN_440 = 5'hd == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_46; 
  wire [4:0] _GEN_441 = 5'he == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_48; 
  wire [4:0] _GEN_442 = 5'hf == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_50; 
  wire [4:0] _GEN_443 = 5'h10 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_52; 
  wire [4:0] _GEN_444 = 5'h11 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_54; 
  wire [4:0] _GEN_445 = 5'h12 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_56; 
  wire [4:0] _GEN_446 = 5'h13 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_58; 
  wire [4:0] _GEN_447 = 5'h14 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_60; 
  wire [4:0] _GEN_448 = 5'h15 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_62; 
  wire [4:0] _GEN_449 = 5'h16 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_64; 
  wire [4:0] _GEN_450 = 5'h17 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_66; 
  wire [4:0] _GEN_451 = 5'h18 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_68; 
  wire [4:0] _GEN_452 = 5'h19 == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_70; 
  wire [4:0] _GEN_453 = 5'h1a == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_72; 
  wire [4:0] _GEN_454 = 5'h1b == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_74; 
  wire [4:0] _GEN_455 = 5'h1c == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_76; 
  wire [4:0] _GEN_456 = 5'h1d == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_78; 
  wire [4:0] _GEN_457 = 5'h1e == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_80; 
  wire [4:0] _GEN_458 = 5'h1f == decoder_if_rd_idx ? _uRegState_io_decoder_if_rd_idx_d_reorder : _GEN_82; 
  wire  _GEN_459 = 5'h0 == decoder_if_rd_idx | _GEN_21; 
  wire  _GEN_460 = 5'h1 == decoder_if_rd_idx | _GEN_23; 
  wire  _GEN_461 = 5'h2 == decoder_if_rd_idx | _GEN_25; 
  wire  _GEN_462 = 5'h3 == decoder_if_rd_idx | _GEN_27; 
  wire  _GEN_463 = 5'h4 == decoder_if_rd_idx | _GEN_29; 
  wire  _GEN_464 = 5'h5 == decoder_if_rd_idx | _GEN_31; 
  wire  _GEN_465 = 5'h6 == decoder_if_rd_idx | _GEN_33; 
  wire  _GEN_466 = 5'h7 == decoder_if_rd_idx | _GEN_35; 
  wire  _GEN_467 = 5'h8 == decoder_if_rd_idx | _GEN_37; 
  wire  _GEN_468 = 5'h9 == decoder_if_rd_idx | _GEN_39; 
  wire  _GEN_469 = 5'ha == decoder_if_rd_idx | _GEN_41; 
  wire  _GEN_470 = 5'hb == decoder_if_rd_idx | _GEN_43; 
  wire  _GEN_471 = 5'hc == decoder_if_rd_idx | _GEN_45; 
  wire  _GEN_472 = 5'hd == decoder_if_rd_idx | _GEN_47; 
  wire  _GEN_473 = 5'he == decoder_if_rd_idx | _GEN_49; 
  wire  _GEN_474 = 5'hf == decoder_if_rd_idx | _GEN_51; 
  wire  _GEN_475 = 5'h10 == decoder_if_rd_idx | _GEN_53; 
  wire  _GEN_476 = 5'h11 == decoder_if_rd_idx | _GEN_55; 
  wire  _GEN_477 = 5'h12 == decoder_if_rd_idx | _GEN_57; 
  wire  _GEN_478 = 5'h13 == decoder_if_rd_idx | _GEN_59; 
  wire  _GEN_479 = 5'h14 == decoder_if_rd_idx | _GEN_61; 
  wire  _GEN_480 = 5'h15 == decoder_if_rd_idx | _GEN_63; 
  wire  _GEN_481 = 5'h16 == decoder_if_rd_idx | _GEN_65; 
  wire  _GEN_482 = 5'h17 == decoder_if_rd_idx | _GEN_67; 
  wire  _GEN_483 = 5'h18 == decoder_if_rd_idx | _GEN_69; 
  wire  _GEN_484 = 5'h19 == decoder_if_rd_idx | _GEN_71; 
  wire  _GEN_485 = 5'h1a == decoder_if_rd_idx | _GEN_73; 
  wire  _GEN_486 = 5'h1b == decoder_if_rd_idx | _GEN_75; 
  wire  _GEN_487 = 5'h1c == decoder_if_rd_idx | _GEN_77; 
  wire  _GEN_488 = 5'h1d == decoder_if_rd_idx | _GEN_79; 
  wire  _GEN_489 = 5'h1e == decoder_if_rd_idx | _GEN_81; 
  wire  _GEN_490 = 5'h1f == decoder_if_rd_idx | _GEN_83; 
  wire [4:0] _GEN_501 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_427 : _GEN_20; 
  wire [4:0] _GEN_502 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_428 : _GEN_22; 
  wire [4:0] _GEN_503 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_429 : _GEN_24; 
  wire [4:0] _GEN_504 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_430 : _GEN_26; 
  wire [4:0] _GEN_505 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_431 : _GEN_28; 
  wire [4:0] _GEN_506 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_432 : _GEN_30; 
  wire [4:0] _GEN_507 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_433 : _GEN_32; 
  wire [4:0] _GEN_508 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_434 : _GEN_34; 
  wire [4:0] _GEN_509 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_435 : _GEN_36; 
  wire [4:0] _GEN_510 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_436 : _GEN_38; 
  wire [4:0] _GEN_511 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_437 : _GEN_40; 
  wire [4:0] _GEN_512 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_438 : _GEN_42; 
  wire [4:0] _GEN_513 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_439 : _GEN_44; 
  wire [4:0] _GEN_514 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_440 : _GEN_46; 
  wire [4:0] _GEN_515 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_441 : _GEN_48; 
  wire [4:0] _GEN_516 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_442 : _GEN_50; 
  wire [4:0] _GEN_517 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_443 : _GEN_52; 
  wire [4:0] _GEN_518 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_444 : _GEN_54; 
  wire [4:0] _GEN_519 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_445 : _GEN_56; 
  wire [4:0] _GEN_520 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_446 : _GEN_58; 
  wire [4:0] _GEN_521 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_447 : _GEN_60; 
  wire [4:0] _GEN_522 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_448 : _GEN_62; 
  wire [4:0] _GEN_523 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_449 : _GEN_64; 
  wire [4:0] _GEN_524 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_450 : _GEN_66; 
  wire [4:0] _GEN_525 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_451 : _GEN_68; 
  wire [4:0] _GEN_526 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_452 : _GEN_70; 
  wire [4:0] _GEN_527 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_453 : _GEN_72; 
  wire [4:0] _GEN_528 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_454 : _GEN_74; 
  wire [4:0] _GEN_529 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_455 : _GEN_76; 
  wire [4:0] _GEN_530 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_456 : _GEN_78; 
  wire [4:0] _GEN_531 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_457 : _GEN_80; 
  wire [4:0] _GEN_532 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_458 : _GEN_82; 
  wire  _GEN_533 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_459 : _GEN_21; 
  wire  _GEN_534 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_460 : _GEN_23; 
  wire  _GEN_535 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_461 : _GEN_25; 
  wire  _GEN_536 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_462 : _GEN_27; 
  wire  _GEN_537 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_463 : _GEN_29; 
  wire  _GEN_538 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_464 : _GEN_31; 
  wire  _GEN_539 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_465 : _GEN_33; 
  wire  _GEN_540 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_466 : _GEN_35; 
  wire  _GEN_541 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_467 : _GEN_37; 
  wire  _GEN_542 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_468 : _GEN_39; 
  wire  _GEN_543 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_469 : _GEN_41; 
  wire  _GEN_544 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_470 : _GEN_43; 
  wire  _GEN_545 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_471 : _GEN_45; 
  wire  _GEN_546 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_472 : _GEN_47; 
  wire  _GEN_547 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_473 : _GEN_49; 
  wire  _GEN_548 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_474 : _GEN_51; 
  wire  _GEN_549 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_475 : _GEN_53; 
  wire  _GEN_550 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_476 : _GEN_55; 
  wire  _GEN_551 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_477 : _GEN_57; 
  wire  _GEN_552 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_478 : _GEN_59; 
  wire  _GEN_553 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_479 : _GEN_61; 
  wire  _GEN_554 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_480 : _GEN_63; 
  wire  _GEN_555 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_481 : _GEN_65; 
  wire  _GEN_556 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_482 : _GEN_67; 
  wire  _GEN_557 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_483 : _GEN_69; 
  wire  _GEN_558 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_484 : _GEN_71; 
  wire  _GEN_559 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_485 : _GEN_73; 
  wire  _GEN_560 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_486 : _GEN_75; 
  wire  _GEN_561 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_487 : _GEN_77; 
  wire  _GEN_562 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_488 : _GEN_79; 
  wire  _GEN_563 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_489 : _GEN_81; 
  wire  _GEN_564 = ~uIntergerRS__io_full & ~uROB__io_full ? _GEN_490 : _GEN_83; 
  wire [4:0] _GEN_1543 = _T_384 ? _GEN_427 : _GEN_20; 
  wire [4:0] _GEN_1544 = _T_384 ? _GEN_428 : _GEN_22; 
  wire [4:0] _GEN_1545 = _T_384 ? _GEN_429 : _GEN_24; 
  wire [4:0] _GEN_1546 = _T_384 ? _GEN_430 : _GEN_26; 
  wire [4:0] _GEN_1547 = _T_384 ? _GEN_431 : _GEN_28; 
  wire [4:0] _GEN_1548 = _T_384 ? _GEN_432 : _GEN_30; 
  wire [4:0] _GEN_1549 = _T_384 ? _GEN_433 : _GEN_32; 
  wire [4:0] _GEN_1550 = _T_384 ? _GEN_434 : _GEN_34; 
  wire [4:0] _GEN_1551 = _T_384 ? _GEN_435 : _GEN_36; 
  wire [4:0] _GEN_1552 = _T_384 ? _GEN_436 : _GEN_38; 
  wire [4:0] _GEN_1553 = _T_384 ? _GEN_437 : _GEN_40; 
  wire [4:0] _GEN_1554 = _T_384 ? _GEN_438 : _GEN_42; 
  wire [4:0] _GEN_1555 = _T_384 ? _GEN_439 : _GEN_44; 
  wire [4:0] _GEN_1556 = _T_384 ? _GEN_440 : _GEN_46; 
  wire [4:0] _GEN_1557 = _T_384 ? _GEN_441 : _GEN_48; 
  wire [4:0] _GEN_1558 = _T_384 ? _GEN_442 : _GEN_50; 
  wire [4:0] _GEN_1559 = _T_384 ? _GEN_443 : _GEN_52; 
  wire [4:0] _GEN_1560 = _T_384 ? _GEN_444 : _GEN_54; 
  wire [4:0] _GEN_1561 = _T_384 ? _GEN_445 : _GEN_56; 
  wire [4:0] _GEN_1562 = _T_384 ? _GEN_446 : _GEN_58; 
  wire [4:0] _GEN_1563 = _T_384 ? _GEN_447 : _GEN_60; 
  wire [4:0] _GEN_1564 = _T_384 ? _GEN_448 : _GEN_62; 
  wire [4:0] _GEN_1565 = _T_384 ? _GEN_449 : _GEN_64; 
  wire [4:0] _GEN_1566 = _T_384 ? _GEN_450 : _GEN_66; 
  wire [4:0] _GEN_1567 = _T_384 ? _GEN_451 : _GEN_68; 
  wire [4:0] _GEN_1568 = _T_384 ? _GEN_452 : _GEN_70; 
  wire [4:0] _GEN_1569 = _T_384 ? _GEN_453 : _GEN_72; 
  wire [4:0] _GEN_1570 = _T_384 ? _GEN_454 : _GEN_74; 
  wire [4:0] _GEN_1571 = _T_384 ? _GEN_455 : _GEN_76; 
  wire [4:0] _GEN_1572 = _T_384 ? _GEN_456 : _GEN_78; 
  wire [4:0] _GEN_1573 = _T_384 ? _GEN_457 : _GEN_80; 
  wire [4:0] _GEN_1574 = _T_384 ? _GEN_458 : _GEN_82; 
  wire  _GEN_1575 = _T_384 ? _GEN_459 : _GEN_21; 
  wire  _GEN_1576 = _T_384 ? _GEN_460 : _GEN_23; 
  wire  _GEN_1577 = _T_384 ? _GEN_461 : _GEN_25; 
  wire  _GEN_1578 = _T_384 ? _GEN_462 : _GEN_27; 
  wire  _GEN_1579 = _T_384 ? _GEN_463 : _GEN_29; 
  wire  _GEN_1580 = _T_384 ? _GEN_464 : _GEN_31; 
  wire  _GEN_1581 = _T_384 ? _GEN_465 : _GEN_33; 
  wire  _GEN_1582 = _T_384 ? _GEN_466 : _GEN_35; 
  wire  _GEN_1583 = _T_384 ? _GEN_467 : _GEN_37; 
  wire  _GEN_1584 = _T_384 ? _GEN_468 : _GEN_39; 
  wire  _GEN_1585 = _T_384 ? _GEN_469 : _GEN_41; 
  wire  _GEN_1586 = _T_384 ? _GEN_470 : _GEN_43; 
  wire  _GEN_1587 = _T_384 ? _GEN_471 : _GEN_45; 
  wire  _GEN_1588 = _T_384 ? _GEN_472 : _GEN_47; 
  wire  _GEN_1589 = _T_384 ? _GEN_473 : _GEN_49; 
  wire  _GEN_1590 = _T_384 ? _GEN_474 : _GEN_51; 
  wire  _GEN_1591 = _T_384 ? _GEN_475 : _GEN_53; 
  wire  _GEN_1592 = _T_384 ? _GEN_476 : _GEN_55; 
  wire  _GEN_1593 = _T_384 ? _GEN_477 : _GEN_57; 
  wire  _GEN_1594 = _T_384 ? _GEN_478 : _GEN_59; 
  wire  _GEN_1595 = _T_384 ? _GEN_479 : _GEN_61; 
  wire  _GEN_1596 = _T_384 ? _GEN_480 : _GEN_63; 
  wire  _GEN_1597 = _T_384 ? _GEN_481 : _GEN_65; 
  wire  _GEN_1598 = _T_384 ? _GEN_482 : _GEN_67; 
  wire  _GEN_1599 = _T_384 ? _GEN_483 : _GEN_69; 
  wire  _GEN_1600 = _T_384 ? _GEN_484 : _GEN_71; 
  wire  _GEN_1601 = _T_384 ? _GEN_485 : _GEN_73; 
  wire  _GEN_1602 = _T_384 ? _GEN_486 : _GEN_75; 
  wire  _GEN_1603 = _T_384 ? _GEN_487 : _GEN_77; 
  wire  _GEN_1604 = _T_384 ? _GEN_488 : _GEN_79; 
  wire  _GEN_1605 = _T_384 ? _GEN_489 : _GEN_81; 
  wire  _GEN_1606 = _T_384 ? _GEN_490 : _GEN_83; 
  wire [4:0] _GEN_2021 = ~uMulDivRS__io_full & _T_351 ? _GEN_427 : _GEN_20; 
  wire [4:0] _GEN_2022 = ~uMulDivRS__io_full & _T_351 ? _GEN_428 : _GEN_22; 
  wire [4:0] _GEN_2023 = ~uMulDivRS__io_full & _T_351 ? _GEN_429 : _GEN_24; 
  wire [4:0] _GEN_2024 = ~uMulDivRS__io_full & _T_351 ? _GEN_430 : _GEN_26; 
  wire [4:0] _GEN_2025 = ~uMulDivRS__io_full & _T_351 ? _GEN_431 : _GEN_28; 
  wire [4:0] _GEN_2026 = ~uMulDivRS__io_full & _T_351 ? _GEN_432 : _GEN_30; 
  wire [4:0] _GEN_2027 = ~uMulDivRS__io_full & _T_351 ? _GEN_433 : _GEN_32; 
  wire [4:0] _GEN_2028 = ~uMulDivRS__io_full & _T_351 ? _GEN_434 : _GEN_34; 
  wire [4:0] _GEN_2029 = ~uMulDivRS__io_full & _T_351 ? _GEN_435 : _GEN_36; 
  wire [4:0] _GEN_2030 = ~uMulDivRS__io_full & _T_351 ? _GEN_436 : _GEN_38; 
  wire [4:0] _GEN_2031 = ~uMulDivRS__io_full & _T_351 ? _GEN_437 : _GEN_40; 
  wire [4:0] _GEN_2032 = ~uMulDivRS__io_full & _T_351 ? _GEN_438 : _GEN_42; 
  wire [4:0] _GEN_2033 = ~uMulDivRS__io_full & _T_351 ? _GEN_439 : _GEN_44; 
  wire [4:0] _GEN_2034 = ~uMulDivRS__io_full & _T_351 ? _GEN_440 : _GEN_46; 
  wire [4:0] _GEN_2035 = ~uMulDivRS__io_full & _T_351 ? _GEN_441 : _GEN_48; 
  wire [4:0] _GEN_2036 = ~uMulDivRS__io_full & _T_351 ? _GEN_442 : _GEN_50; 
  wire [4:0] _GEN_2037 = ~uMulDivRS__io_full & _T_351 ? _GEN_443 : _GEN_52; 
  wire [4:0] _GEN_2038 = ~uMulDivRS__io_full & _T_351 ? _GEN_444 : _GEN_54; 
  wire [4:0] _GEN_2039 = ~uMulDivRS__io_full & _T_351 ? _GEN_445 : _GEN_56; 
  wire [4:0] _GEN_2040 = ~uMulDivRS__io_full & _T_351 ? _GEN_446 : _GEN_58; 
  wire [4:0] _GEN_2041 = ~uMulDivRS__io_full & _T_351 ? _GEN_447 : _GEN_60; 
  wire [4:0] _GEN_2042 = ~uMulDivRS__io_full & _T_351 ? _GEN_448 : _GEN_62; 
  wire [4:0] _GEN_2043 = ~uMulDivRS__io_full & _T_351 ? _GEN_449 : _GEN_64; 
  wire [4:0] _GEN_2044 = ~uMulDivRS__io_full & _T_351 ? _GEN_450 : _GEN_66; 
  wire [4:0] _GEN_2045 = ~uMulDivRS__io_full & _T_351 ? _GEN_451 : _GEN_68; 
  wire [4:0] _GEN_2046 = ~uMulDivRS__io_full & _T_351 ? _GEN_452 : _GEN_70; 
  wire [4:0] _GEN_2047 = ~uMulDivRS__io_full & _T_351 ? _GEN_453 : _GEN_72; 
  wire [4:0] _GEN_2048 = ~uMulDivRS__io_full & _T_351 ? _GEN_454 : _GEN_74; 
  wire [4:0] _GEN_2049 = ~uMulDivRS__io_full & _T_351 ? _GEN_455 : _GEN_76; 
  wire [4:0] _GEN_2050 = ~uMulDivRS__io_full & _T_351 ? _GEN_456 : _GEN_78; 
  wire [4:0] _GEN_2051 = ~uMulDivRS__io_full & _T_351 ? _GEN_457 : _GEN_80; 
  wire [4:0] _GEN_2052 = ~uMulDivRS__io_full & _T_351 ? _GEN_458 : _GEN_82; 
  wire  _GEN_2053 = ~uMulDivRS__io_full & _T_351 ? _GEN_459 : _GEN_21; 
  wire  _GEN_2054 = ~uMulDivRS__io_full & _T_351 ? _GEN_460 : _GEN_23; 
  wire  _GEN_2055 = ~uMulDivRS__io_full & _T_351 ? _GEN_461 : _GEN_25; 
  wire  _GEN_2056 = ~uMulDivRS__io_full & _T_351 ? _GEN_462 : _GEN_27; 
  wire  _GEN_2057 = ~uMulDivRS__io_full & _T_351 ? _GEN_463 : _GEN_29; 
  wire  _GEN_2058 = ~uMulDivRS__io_full & _T_351 ? _GEN_464 : _GEN_31; 
  wire  _GEN_2059 = ~uMulDivRS__io_full & _T_351 ? _GEN_465 : _GEN_33; 
  wire  _GEN_2060 = ~uMulDivRS__io_full & _T_351 ? _GEN_466 : _GEN_35; 
  wire  _GEN_2061 = ~uMulDivRS__io_full & _T_351 ? _GEN_467 : _GEN_37; 
  wire  _GEN_2062 = ~uMulDivRS__io_full & _T_351 ? _GEN_468 : _GEN_39; 
  wire  _GEN_2063 = ~uMulDivRS__io_full & _T_351 ? _GEN_469 : _GEN_41; 
  wire  _GEN_2064 = ~uMulDivRS__io_full & _T_351 ? _GEN_470 : _GEN_43; 
  wire  _GEN_2065 = ~uMulDivRS__io_full & _T_351 ? _GEN_471 : _GEN_45; 
  wire  _GEN_2066 = ~uMulDivRS__io_full & _T_351 ? _GEN_472 : _GEN_47; 
  wire  _GEN_2067 = ~uMulDivRS__io_full & _T_351 ? _GEN_473 : _GEN_49; 
  wire  _GEN_2068 = ~uMulDivRS__io_full & _T_351 ? _GEN_474 : _GEN_51; 
  wire  _GEN_2069 = ~uMulDivRS__io_full & _T_351 ? _GEN_475 : _GEN_53; 
  wire  _GEN_2070 = ~uMulDivRS__io_full & _T_351 ? _GEN_476 : _GEN_55; 
  wire  _GEN_2071 = ~uMulDivRS__io_full & _T_351 ? _GEN_477 : _GEN_57; 
  wire  _GEN_2072 = ~uMulDivRS__io_full & _T_351 ? _GEN_478 : _GEN_59; 
  wire  _GEN_2073 = ~uMulDivRS__io_full & _T_351 ? _GEN_479 : _GEN_61; 
  wire  _GEN_2074 = ~uMulDivRS__io_full & _T_351 ? _GEN_480 : _GEN_63; 
  wire  _GEN_2075 = ~uMulDivRS__io_full & _T_351 ? _GEN_481 : _GEN_65; 
  wire  _GEN_2076 = ~uMulDivRS__io_full & _T_351 ? _GEN_482 : _GEN_67; 
  wire  _GEN_2077 = ~uMulDivRS__io_full & _T_351 ? _GEN_483 : _GEN_69; 
  wire  _GEN_2078 = ~uMulDivRS__io_full & _T_351 ? _GEN_484 : _GEN_71; 
  wire  _GEN_2079 = ~uMulDivRS__io_full & _T_351 ? _GEN_485 : _GEN_73; 
  wire  _GEN_2080 = ~uMulDivRS__io_full & _T_351 ? _GEN_486 : _GEN_75; 
  wire  _GEN_2081 = ~uMulDivRS__io_full & _T_351 ? _GEN_487 : _GEN_77; 
  wire  _GEN_2082 = ~uMulDivRS__io_full & _T_351 ? _GEN_488 : _GEN_79; 
  wire  _GEN_2083 = ~uMulDivRS__io_full & _T_351 ? _GEN_489 : _GEN_81; 
  wire  _GEN_2084 = ~uMulDivRS__io_full & _T_351 ? _GEN_490 : _GEN_83; 
  wire [4:0] _GEN_2095 = muldiv_inst_r_io_d ? _GEN_2021 : _GEN_20; 
  wire [4:0] _GEN_2096 = muldiv_inst_r_io_d ? _GEN_2022 : _GEN_22; 
  wire [4:0] _GEN_2097 = muldiv_inst_r_io_d ? _GEN_2023 : _GEN_24; 
  wire [4:0] _GEN_2098 = muldiv_inst_r_io_d ? _GEN_2024 : _GEN_26; 
  wire [4:0] _GEN_2099 = muldiv_inst_r_io_d ? _GEN_2025 : _GEN_28; 
  wire [4:0] _GEN_2100 = muldiv_inst_r_io_d ? _GEN_2026 : _GEN_30; 
  wire [4:0] _GEN_2101 = muldiv_inst_r_io_d ? _GEN_2027 : _GEN_32; 
  wire [4:0] _GEN_2102 = muldiv_inst_r_io_d ? _GEN_2028 : _GEN_34; 
  wire [4:0] _GEN_2103 = muldiv_inst_r_io_d ? _GEN_2029 : _GEN_36; 
  wire [4:0] _GEN_2104 = muldiv_inst_r_io_d ? _GEN_2030 : _GEN_38; 
  wire [4:0] _GEN_2105 = muldiv_inst_r_io_d ? _GEN_2031 : _GEN_40; 
  wire [4:0] _GEN_2106 = muldiv_inst_r_io_d ? _GEN_2032 : _GEN_42; 
  wire [4:0] _GEN_2107 = muldiv_inst_r_io_d ? _GEN_2033 : _GEN_44; 
  wire [4:0] _GEN_2108 = muldiv_inst_r_io_d ? _GEN_2034 : _GEN_46; 
  wire [4:0] _GEN_2109 = muldiv_inst_r_io_d ? _GEN_2035 : _GEN_48; 
  wire [4:0] _GEN_2110 = muldiv_inst_r_io_d ? _GEN_2036 : _GEN_50; 
  wire [4:0] _GEN_2111 = muldiv_inst_r_io_d ? _GEN_2037 : _GEN_52; 
  wire [4:0] _GEN_2112 = muldiv_inst_r_io_d ? _GEN_2038 : _GEN_54; 
  wire [4:0] _GEN_2113 = muldiv_inst_r_io_d ? _GEN_2039 : _GEN_56; 
  wire [4:0] _GEN_2114 = muldiv_inst_r_io_d ? _GEN_2040 : _GEN_58; 
  wire [4:0] _GEN_2115 = muldiv_inst_r_io_d ? _GEN_2041 : _GEN_60; 
  wire [4:0] _GEN_2116 = muldiv_inst_r_io_d ? _GEN_2042 : _GEN_62; 
  wire [4:0] _GEN_2117 = muldiv_inst_r_io_d ? _GEN_2043 : _GEN_64; 
  wire [4:0] _GEN_2118 = muldiv_inst_r_io_d ? _GEN_2044 : _GEN_66; 
  wire [4:0] _GEN_2119 = muldiv_inst_r_io_d ? _GEN_2045 : _GEN_68; 
  wire [4:0] _GEN_2120 = muldiv_inst_r_io_d ? _GEN_2046 : _GEN_70; 
  wire [4:0] _GEN_2121 = muldiv_inst_r_io_d ? _GEN_2047 : _GEN_72; 
  wire [4:0] _GEN_2122 = muldiv_inst_r_io_d ? _GEN_2048 : _GEN_74; 
  wire [4:0] _GEN_2123 = muldiv_inst_r_io_d ? _GEN_2049 : _GEN_76; 
  wire [4:0] _GEN_2124 = muldiv_inst_r_io_d ? _GEN_2050 : _GEN_78; 
  wire [4:0] _GEN_2125 = muldiv_inst_r_io_d ? _GEN_2051 : _GEN_80; 
  wire [4:0] _GEN_2126 = muldiv_inst_r_io_d ? _GEN_2052 : _GEN_82; 
  wire  _GEN_2127 = muldiv_inst_r_io_d ? _GEN_2053 : _GEN_21; 
  wire  _GEN_2128 = muldiv_inst_r_io_d ? _GEN_2054 : _GEN_23; 
  wire  _GEN_2129 = muldiv_inst_r_io_d ? _GEN_2055 : _GEN_25; 
  wire  _GEN_2130 = muldiv_inst_r_io_d ? _GEN_2056 : _GEN_27; 
  wire  _GEN_2131 = muldiv_inst_r_io_d ? _GEN_2057 : _GEN_29; 
  wire  _GEN_2132 = muldiv_inst_r_io_d ? _GEN_2058 : _GEN_31; 
  wire  _GEN_2133 = muldiv_inst_r_io_d ? _GEN_2059 : _GEN_33; 
  wire  _GEN_2134 = muldiv_inst_r_io_d ? _GEN_2060 : _GEN_35; 
  wire  _GEN_2135 = muldiv_inst_r_io_d ? _GEN_2061 : _GEN_37; 
  wire  _GEN_2136 = muldiv_inst_r_io_d ? _GEN_2062 : _GEN_39; 
  wire  _GEN_2137 = muldiv_inst_r_io_d ? _GEN_2063 : _GEN_41; 
  wire  _GEN_2138 = muldiv_inst_r_io_d ? _GEN_2064 : _GEN_43; 
  wire  _GEN_2139 = muldiv_inst_r_io_d ? _GEN_2065 : _GEN_45; 
  wire  _GEN_2140 = muldiv_inst_r_io_d ? _GEN_2066 : _GEN_47; 
  wire  _GEN_2141 = muldiv_inst_r_io_d ? _GEN_2067 : _GEN_49; 
  wire  _GEN_2142 = muldiv_inst_r_io_d ? _GEN_2068 : _GEN_51; 
  wire  _GEN_2143 = muldiv_inst_r_io_d ? _GEN_2069 : _GEN_53; 
  wire  _GEN_2144 = muldiv_inst_r_io_d ? _GEN_2070 : _GEN_55; 
  wire  _GEN_2145 = muldiv_inst_r_io_d ? _GEN_2071 : _GEN_57; 
  wire  _GEN_2146 = muldiv_inst_r_io_d ? _GEN_2072 : _GEN_59; 
  wire  _GEN_2147 = muldiv_inst_r_io_d ? _GEN_2073 : _GEN_61; 
  wire  _GEN_2148 = muldiv_inst_r_io_d ? _GEN_2074 : _GEN_63; 
  wire  _GEN_2149 = muldiv_inst_r_io_d ? _GEN_2075 : _GEN_65; 
  wire  _GEN_2150 = muldiv_inst_r_io_d ? _GEN_2076 : _GEN_67; 
  wire  _GEN_2151 = muldiv_inst_r_io_d ? _GEN_2077 : _GEN_69; 
  wire  _GEN_2152 = muldiv_inst_r_io_d ? _GEN_2078 : _GEN_71; 
  wire  _GEN_2153 = muldiv_inst_r_io_d ? _GEN_2079 : _GEN_73; 
  wire  _GEN_2154 = muldiv_inst_r_io_d ? _GEN_2080 : _GEN_75; 
  wire  _GEN_2155 = muldiv_inst_r_io_d ? _GEN_2081 : _GEN_77; 
  wire  _GEN_2156 = muldiv_inst_r_io_d ? _GEN_2082 : _GEN_79; 
  wire  _GEN_2157 = muldiv_inst_r_io_d ? _GEN_2083 : _GEN_81; 
  wire  _GEN_2158 = muldiv_inst_r_io_d ? _GEN_2084 : _GEN_83; 
  wire  _GEN_2159 = load_inst_r_io_d ? _T_384 : _GEN_2085; 
  wire [4:0] _GEN_2171 = load_inst_r_io_d ? _GEN_1543 : _GEN_2095; 
  wire [4:0] _GEN_2172 = load_inst_r_io_d ? _GEN_1544 : _GEN_2096; 
  wire [4:0] _GEN_2173 = load_inst_r_io_d ? _GEN_1545 : _GEN_2097; 
  wire [4:0] _GEN_2174 = load_inst_r_io_d ? _GEN_1546 : _GEN_2098; 
  wire [4:0] _GEN_2175 = load_inst_r_io_d ? _GEN_1547 : _GEN_2099; 
  wire [4:0] _GEN_2176 = load_inst_r_io_d ? _GEN_1548 : _GEN_2100; 
  wire [4:0] _GEN_2177 = load_inst_r_io_d ? _GEN_1549 : _GEN_2101; 
  wire [4:0] _GEN_2178 = load_inst_r_io_d ? _GEN_1550 : _GEN_2102; 
  wire [4:0] _GEN_2179 = load_inst_r_io_d ? _GEN_1551 : _GEN_2103; 
  wire [4:0] _GEN_2180 = load_inst_r_io_d ? _GEN_1552 : _GEN_2104; 
  wire [4:0] _GEN_2181 = load_inst_r_io_d ? _GEN_1553 : _GEN_2105; 
  wire [4:0] _GEN_2182 = load_inst_r_io_d ? _GEN_1554 : _GEN_2106; 
  wire [4:0] _GEN_2183 = load_inst_r_io_d ? _GEN_1555 : _GEN_2107; 
  wire [4:0] _GEN_2184 = load_inst_r_io_d ? _GEN_1556 : _GEN_2108; 
  wire [4:0] _GEN_2185 = load_inst_r_io_d ? _GEN_1557 : _GEN_2109; 
  wire [4:0] _GEN_2186 = load_inst_r_io_d ? _GEN_1558 : _GEN_2110; 
  wire [4:0] _GEN_2187 = load_inst_r_io_d ? _GEN_1559 : _GEN_2111; 
  wire [4:0] _GEN_2188 = load_inst_r_io_d ? _GEN_1560 : _GEN_2112; 
  wire [4:0] _GEN_2189 = load_inst_r_io_d ? _GEN_1561 : _GEN_2113; 
  wire [4:0] _GEN_2190 = load_inst_r_io_d ? _GEN_1562 : _GEN_2114; 
  wire [4:0] _GEN_2191 = load_inst_r_io_d ? _GEN_1563 : _GEN_2115; 
  wire [4:0] _GEN_2192 = load_inst_r_io_d ? _GEN_1564 : _GEN_2116; 
  wire [4:0] _GEN_2193 = load_inst_r_io_d ? _GEN_1565 : _GEN_2117; 
  wire [4:0] _GEN_2194 = load_inst_r_io_d ? _GEN_1566 : _GEN_2118; 
  wire [4:0] _GEN_2195 = load_inst_r_io_d ? _GEN_1567 : _GEN_2119; 
  wire [4:0] _GEN_2196 = load_inst_r_io_d ? _GEN_1568 : _GEN_2120; 
  wire [4:0] _GEN_2197 = load_inst_r_io_d ? _GEN_1569 : _GEN_2121; 
  wire [4:0] _GEN_2198 = load_inst_r_io_d ? _GEN_1570 : _GEN_2122; 
  wire [4:0] _GEN_2199 = load_inst_r_io_d ? _GEN_1571 : _GEN_2123; 
  wire [4:0] _GEN_2200 = load_inst_r_io_d ? _GEN_1572 : _GEN_2124; 
  wire [4:0] _GEN_2201 = load_inst_r_io_d ? _GEN_1573 : _GEN_2125; 
  wire [4:0] _GEN_2202 = load_inst_r_io_d ? _GEN_1574 : _GEN_2126; 
  wire  _GEN_2203 = load_inst_r_io_d ? _GEN_1575 : _GEN_2127; 
  wire  _GEN_2204 = load_inst_r_io_d ? _GEN_1576 : _GEN_2128; 
  wire  _GEN_2205 = load_inst_r_io_d ? _GEN_1577 : _GEN_2129; 
  wire  _GEN_2206 = load_inst_r_io_d ? _GEN_1578 : _GEN_2130; 
  wire  _GEN_2207 = load_inst_r_io_d ? _GEN_1579 : _GEN_2131; 
  wire  _GEN_2208 = load_inst_r_io_d ? _GEN_1580 : _GEN_2132; 
  wire  _GEN_2209 = load_inst_r_io_d ? _GEN_1581 : _GEN_2133; 
  wire  _GEN_2210 = load_inst_r_io_d ? _GEN_1582 : _GEN_2134; 
  wire  _GEN_2211 = load_inst_r_io_d ? _GEN_1583 : _GEN_2135; 
  wire  _GEN_2212 = load_inst_r_io_d ? _GEN_1584 : _GEN_2136; 
  wire  _GEN_2213 = load_inst_r_io_d ? _GEN_1585 : _GEN_2137; 
  wire  _GEN_2214 = load_inst_r_io_d ? _GEN_1586 : _GEN_2138; 
  wire  _GEN_2215 = load_inst_r_io_d ? _GEN_1587 : _GEN_2139; 
  wire  _GEN_2216 = load_inst_r_io_d ? _GEN_1588 : _GEN_2140; 
  wire  _GEN_2217 = load_inst_r_io_d ? _GEN_1589 : _GEN_2141; 
  wire  _GEN_2218 = load_inst_r_io_d ? _GEN_1590 : _GEN_2142; 
  wire  _GEN_2219 = load_inst_r_io_d ? _GEN_1591 : _GEN_2143; 
  wire  _GEN_2220 = load_inst_r_io_d ? _GEN_1592 : _GEN_2144; 
  wire  _GEN_2221 = load_inst_r_io_d ? _GEN_1593 : _GEN_2145; 
  wire  _GEN_2222 = load_inst_r_io_d ? _GEN_1594 : _GEN_2146; 
  wire  _GEN_2223 = load_inst_r_io_d ? _GEN_1595 : _GEN_2147; 
  wire  _GEN_2224 = load_inst_r_io_d ? _GEN_1596 : _GEN_2148; 
  wire  _GEN_2225 = load_inst_r_io_d ? _GEN_1597 : _GEN_2149; 
  wire  _GEN_2226 = load_inst_r_io_d ? _GEN_1598 : _GEN_2150; 
  wire  _GEN_2227 = load_inst_r_io_d ? _GEN_1599 : _GEN_2151; 
  wire  _GEN_2228 = load_inst_r_io_d ? _GEN_1600 : _GEN_2152; 
  wire  _GEN_2229 = load_inst_r_io_d ? _GEN_1601 : _GEN_2153; 
  wire  _GEN_2230 = load_inst_r_io_d ? _GEN_1602 : _GEN_2154; 
  wire  _GEN_2231 = load_inst_r_io_d ? _GEN_1603 : _GEN_2155; 
  wire  _GEN_2232 = load_inst_r_io_d ? _GEN_1604 : _GEN_2156; 
  wire  _GEN_2233 = load_inst_r_io_d ? _GEN_1605 : _GEN_2157; 
  wire  _GEN_2234 = load_inst_r_io_d ? _GEN_1606 : _GEN_2158; 
  wire  _GEN_2242 = store_inst_r_io_d ? _T_384 : _GEN_2159; 
  wire [4:0] _GEN_2254 = store_inst_r_io_d ? _GEN_20 : _GEN_2171; 
  wire [4:0] _GEN_2255 = store_inst_r_io_d ? _GEN_22 : _GEN_2172; 
  wire [4:0] _GEN_2256 = store_inst_r_io_d ? _GEN_24 : _GEN_2173; 
  wire [4:0] _GEN_2257 = store_inst_r_io_d ? _GEN_26 : _GEN_2174; 
  wire [4:0] _GEN_2258 = store_inst_r_io_d ? _GEN_28 : _GEN_2175; 
  wire [4:0] _GEN_2259 = store_inst_r_io_d ? _GEN_30 : _GEN_2176; 
  wire [4:0] _GEN_2260 = store_inst_r_io_d ? _GEN_32 : _GEN_2177; 
  wire [4:0] _GEN_2261 = store_inst_r_io_d ? _GEN_34 : _GEN_2178; 
  wire [4:0] _GEN_2262 = store_inst_r_io_d ? _GEN_36 : _GEN_2179; 
  wire [4:0] _GEN_2263 = store_inst_r_io_d ? _GEN_38 : _GEN_2180; 
  wire [4:0] _GEN_2264 = store_inst_r_io_d ? _GEN_40 : _GEN_2181; 
  wire [4:0] _GEN_2265 = store_inst_r_io_d ? _GEN_42 : _GEN_2182; 
  wire [4:0] _GEN_2266 = store_inst_r_io_d ? _GEN_44 : _GEN_2183; 
  wire [4:0] _GEN_2267 = store_inst_r_io_d ? _GEN_46 : _GEN_2184; 
  wire [4:0] _GEN_2268 = store_inst_r_io_d ? _GEN_48 : _GEN_2185; 
  wire [4:0] _GEN_2269 = store_inst_r_io_d ? _GEN_50 : _GEN_2186; 
  wire [4:0] _GEN_2270 = store_inst_r_io_d ? _GEN_52 : _GEN_2187; 
  wire [4:0] _GEN_2271 = store_inst_r_io_d ? _GEN_54 : _GEN_2188; 
  wire [4:0] _GEN_2272 = store_inst_r_io_d ? _GEN_56 : _GEN_2189; 
  wire [4:0] _GEN_2273 = store_inst_r_io_d ? _GEN_58 : _GEN_2190; 
  wire [4:0] _GEN_2274 = store_inst_r_io_d ? _GEN_60 : _GEN_2191; 
  wire [4:0] _GEN_2275 = store_inst_r_io_d ? _GEN_62 : _GEN_2192; 
  wire [4:0] _GEN_2276 = store_inst_r_io_d ? _GEN_64 : _GEN_2193; 
  wire [4:0] _GEN_2277 = store_inst_r_io_d ? _GEN_66 : _GEN_2194; 
  wire [4:0] _GEN_2278 = store_inst_r_io_d ? _GEN_68 : _GEN_2195; 
  wire [4:0] _GEN_2279 = store_inst_r_io_d ? _GEN_70 : _GEN_2196; 
  wire [4:0] _GEN_2280 = store_inst_r_io_d ? _GEN_72 : _GEN_2197; 
  wire [4:0] _GEN_2281 = store_inst_r_io_d ? _GEN_74 : _GEN_2198; 
  wire [4:0] _GEN_2282 = store_inst_r_io_d ? _GEN_76 : _GEN_2199; 
  wire [4:0] _GEN_2283 = store_inst_r_io_d ? _GEN_78 : _GEN_2200; 
  wire [4:0] _GEN_2284 = store_inst_r_io_d ? _GEN_80 : _GEN_2201; 
  wire [4:0] _GEN_2285 = store_inst_r_io_d ? _GEN_82 : _GEN_2202; 
  wire  _GEN_2286 = store_inst_r_io_d ? _GEN_21 : _GEN_2203; 
  wire  _GEN_2287 = store_inst_r_io_d ? _GEN_23 : _GEN_2204; 
  wire  _GEN_2288 = store_inst_r_io_d ? _GEN_25 : _GEN_2205; 
  wire  _GEN_2289 = store_inst_r_io_d ? _GEN_27 : _GEN_2206; 
  wire  _GEN_2290 = store_inst_r_io_d ? _GEN_29 : _GEN_2207; 
  wire  _GEN_2291 = store_inst_r_io_d ? _GEN_31 : _GEN_2208; 
  wire  _GEN_2292 = store_inst_r_io_d ? _GEN_33 : _GEN_2209; 
  wire  _GEN_2293 = store_inst_r_io_d ? _GEN_35 : _GEN_2210; 
  wire  _GEN_2294 = store_inst_r_io_d ? _GEN_37 : _GEN_2211; 
  wire  _GEN_2295 = store_inst_r_io_d ? _GEN_39 : _GEN_2212; 
  wire  _GEN_2296 = store_inst_r_io_d ? _GEN_41 : _GEN_2213; 
  wire  _GEN_2297 = store_inst_r_io_d ? _GEN_43 : _GEN_2214; 
  wire  _GEN_2298 = store_inst_r_io_d ? _GEN_45 : _GEN_2215; 
  wire  _GEN_2299 = store_inst_r_io_d ? _GEN_47 : _GEN_2216; 
  wire  _GEN_2300 = store_inst_r_io_d ? _GEN_49 : _GEN_2217; 
  wire  _GEN_2301 = store_inst_r_io_d ? _GEN_51 : _GEN_2218; 
  wire  _GEN_2302 = store_inst_r_io_d ? _GEN_53 : _GEN_2219; 
  wire  _GEN_2303 = store_inst_r_io_d ? _GEN_55 : _GEN_2220; 
  wire  _GEN_2304 = store_inst_r_io_d ? _GEN_57 : _GEN_2221; 
  wire  _GEN_2305 = store_inst_r_io_d ? _GEN_59 : _GEN_2222; 
  wire  _GEN_2306 = store_inst_r_io_d ? _GEN_61 : _GEN_2223; 
  wire  _GEN_2307 = store_inst_r_io_d ? _GEN_63 : _GEN_2224; 
  wire  _GEN_2308 = store_inst_r_io_d ? _GEN_65 : _GEN_2225; 
  wire  _GEN_2309 = store_inst_r_io_d ? _GEN_67 : _GEN_2226; 
  wire  _GEN_2310 = store_inst_r_io_d ? _GEN_69 : _GEN_2227; 
  wire  _GEN_2311 = store_inst_r_io_d ? _GEN_71 : _GEN_2228; 
  wire  _GEN_2312 = store_inst_r_io_d ? _GEN_73 : _GEN_2229; 
  wire  _GEN_2313 = store_inst_r_io_d ? _GEN_75 : _GEN_2230; 
  wire  _GEN_2314 = store_inst_r_io_d ? _GEN_77 : _GEN_2231; 
  wire  _GEN_2315 = store_inst_r_io_d ? _GEN_79 : _GEN_2232; 
  wire  _GEN_2316 = store_inst_r_io_d ? _GEN_81 : _GEN_2233; 
  wire  _GEN_2317 = store_inst_r_io_d ? _GEN_83 : _GEN_2234; 
  wire  _GEN_2325 = branch_inst_r_io_d ? _T_352 : _GEN_2242; 
  wire [4:0] _GEN_2344 = branch_inst_r_io_d ? _GEN_20 : _GEN_2254; 
  wire [4:0] _GEN_2345 = branch_inst_r_io_d ? _GEN_22 : _GEN_2255; 
  wire [4:0] _GEN_2346 = branch_inst_r_io_d ? _GEN_24 : _GEN_2256; 
  wire [4:0] _GEN_2347 = branch_inst_r_io_d ? _GEN_26 : _GEN_2257; 
  wire [4:0] _GEN_2348 = branch_inst_r_io_d ? _GEN_28 : _GEN_2258; 
  wire [4:0] _GEN_2349 = branch_inst_r_io_d ? _GEN_30 : _GEN_2259; 
  wire [4:0] _GEN_2350 = branch_inst_r_io_d ? _GEN_32 : _GEN_2260; 
  wire [4:0] _GEN_2351 = branch_inst_r_io_d ? _GEN_34 : _GEN_2261; 
  wire [4:0] _GEN_2352 = branch_inst_r_io_d ? _GEN_36 : _GEN_2262; 
  wire [4:0] _GEN_2353 = branch_inst_r_io_d ? _GEN_38 : _GEN_2263; 
  wire [4:0] _GEN_2354 = branch_inst_r_io_d ? _GEN_40 : _GEN_2264; 
  wire [4:0] _GEN_2355 = branch_inst_r_io_d ? _GEN_42 : _GEN_2265; 
  wire [4:0] _GEN_2356 = branch_inst_r_io_d ? _GEN_44 : _GEN_2266; 
  wire [4:0] _GEN_2357 = branch_inst_r_io_d ? _GEN_46 : _GEN_2267; 
  wire [4:0] _GEN_2358 = branch_inst_r_io_d ? _GEN_48 : _GEN_2268; 
  wire [4:0] _GEN_2359 = branch_inst_r_io_d ? _GEN_50 : _GEN_2269; 
  wire [4:0] _GEN_2360 = branch_inst_r_io_d ? _GEN_52 : _GEN_2270; 
  wire [4:0] _GEN_2361 = branch_inst_r_io_d ? _GEN_54 : _GEN_2271; 
  wire [4:0] _GEN_2362 = branch_inst_r_io_d ? _GEN_56 : _GEN_2272; 
  wire [4:0] _GEN_2363 = branch_inst_r_io_d ? _GEN_58 : _GEN_2273; 
  wire [4:0] _GEN_2364 = branch_inst_r_io_d ? _GEN_60 : _GEN_2274; 
  wire [4:0] _GEN_2365 = branch_inst_r_io_d ? _GEN_62 : _GEN_2275; 
  wire [4:0] _GEN_2366 = branch_inst_r_io_d ? _GEN_64 : _GEN_2276; 
  wire [4:0] _GEN_2367 = branch_inst_r_io_d ? _GEN_66 : _GEN_2277; 
  wire [4:0] _GEN_2368 = branch_inst_r_io_d ? _GEN_68 : _GEN_2278; 
  wire [4:0] _GEN_2369 = branch_inst_r_io_d ? _GEN_70 : _GEN_2279; 
  wire [4:0] _GEN_2370 = branch_inst_r_io_d ? _GEN_72 : _GEN_2280; 
  wire [4:0] _GEN_2371 = branch_inst_r_io_d ? _GEN_74 : _GEN_2281; 
  wire [4:0] _GEN_2372 = branch_inst_r_io_d ? _GEN_76 : _GEN_2282; 
  wire [4:0] _GEN_2373 = branch_inst_r_io_d ? _GEN_78 : _GEN_2283; 
  wire [4:0] _GEN_2374 = branch_inst_r_io_d ? _GEN_80 : _GEN_2284; 
  wire [4:0] _GEN_2375 = branch_inst_r_io_d ? _GEN_82 : _GEN_2285; 
  wire  _GEN_2376 = branch_inst_r_io_d ? _GEN_21 : _GEN_2286; 
  wire  _GEN_2377 = branch_inst_r_io_d ? _GEN_23 : _GEN_2287; 
  wire  _GEN_2378 = branch_inst_r_io_d ? _GEN_25 : _GEN_2288; 
  wire  _GEN_2379 = branch_inst_r_io_d ? _GEN_27 : _GEN_2289; 
  wire  _GEN_2380 = branch_inst_r_io_d ? _GEN_29 : _GEN_2290; 
  wire  _GEN_2381 = branch_inst_r_io_d ? _GEN_31 : _GEN_2291; 
  wire  _GEN_2382 = branch_inst_r_io_d ? _GEN_33 : _GEN_2292; 
  wire  _GEN_2383 = branch_inst_r_io_d ? _GEN_35 : _GEN_2293; 
  wire  _GEN_2384 = branch_inst_r_io_d ? _GEN_37 : _GEN_2294; 
  wire  _GEN_2385 = branch_inst_r_io_d ? _GEN_39 : _GEN_2295; 
  wire  _GEN_2386 = branch_inst_r_io_d ? _GEN_41 : _GEN_2296; 
  wire  _GEN_2387 = branch_inst_r_io_d ? _GEN_43 : _GEN_2297; 
  wire  _GEN_2388 = branch_inst_r_io_d ? _GEN_45 : _GEN_2298; 
  wire  _GEN_2389 = branch_inst_r_io_d ? _GEN_47 : _GEN_2299; 
  wire  _GEN_2390 = branch_inst_r_io_d ? _GEN_49 : _GEN_2300; 
  wire  _GEN_2391 = branch_inst_r_io_d ? _GEN_51 : _GEN_2301; 
  wire  _GEN_2392 = branch_inst_r_io_d ? _GEN_53 : _GEN_2302; 
  wire  _GEN_2393 = branch_inst_r_io_d ? _GEN_55 : _GEN_2303; 
  wire  _GEN_2394 = branch_inst_r_io_d ? _GEN_57 : _GEN_2304; 
  wire  _GEN_2395 = branch_inst_r_io_d ? _GEN_59 : _GEN_2305; 
  wire  _GEN_2396 = branch_inst_r_io_d ? _GEN_61 : _GEN_2306; 
  wire  _GEN_2397 = branch_inst_r_io_d ? _GEN_63 : _GEN_2307; 
  wire  _GEN_2398 = branch_inst_r_io_d ? _GEN_65 : _GEN_2308; 
  wire  _GEN_2399 = branch_inst_r_io_d ? _GEN_67 : _GEN_2309; 
  wire  _GEN_2400 = branch_inst_r_io_d ? _GEN_69 : _GEN_2310; 
  wire  _GEN_2401 = branch_inst_r_io_d ? _GEN_71 : _GEN_2311; 
  wire  _GEN_2402 = branch_inst_r_io_d ? _GEN_73 : _GEN_2312; 
  wire  _GEN_2403 = branch_inst_r_io_d ? _GEN_75 : _GEN_2313; 
  wire  _GEN_2404 = branch_inst_r_io_d ? _GEN_77 : _GEN_2314; 
  wire  _GEN_2405 = branch_inst_r_io_d ? _GEN_79 : _GEN_2315; 
  wire  _GEN_2406 = branch_inst_r_io_d ? _GEN_81 : _GEN_2316; 
  wire  _GEN_2407 = branch_inst_r_io_d ? _GEN_83 : _GEN_2317; 
  wire  _GEN_2415 = integer_inst_r_io_d ? _T_352 : _GEN_2325; 
  wire [4:0] _GEN_2426 = integer_inst_r_io_d ? _GEN_501 : _GEN_2344; 
  wire [4:0] _GEN_2427 = integer_inst_r_io_d ? _GEN_502 : _GEN_2345; 
  wire [4:0] _GEN_2428 = integer_inst_r_io_d ? _GEN_503 : _GEN_2346; 
  wire [4:0] _GEN_2429 = integer_inst_r_io_d ? _GEN_504 : _GEN_2347; 
  wire [4:0] _GEN_2430 = integer_inst_r_io_d ? _GEN_505 : _GEN_2348; 
  wire [4:0] _GEN_2431 = integer_inst_r_io_d ? _GEN_506 : _GEN_2349; 
  wire [4:0] _GEN_2432 = integer_inst_r_io_d ? _GEN_507 : _GEN_2350; 
  wire [4:0] _GEN_2433 = integer_inst_r_io_d ? _GEN_508 : _GEN_2351; 
  wire [4:0] _GEN_2434 = integer_inst_r_io_d ? _GEN_509 : _GEN_2352; 
  wire [4:0] _GEN_2435 = integer_inst_r_io_d ? _GEN_510 : _GEN_2353; 
  wire [4:0] _GEN_2436 = integer_inst_r_io_d ? _GEN_511 : _GEN_2354; 
  wire [4:0] _GEN_2437 = integer_inst_r_io_d ? _GEN_512 : _GEN_2355; 
  wire [4:0] _GEN_2438 = integer_inst_r_io_d ? _GEN_513 : _GEN_2356; 
  wire [4:0] _GEN_2439 = integer_inst_r_io_d ? _GEN_514 : _GEN_2357; 
  wire [4:0] _GEN_2440 = integer_inst_r_io_d ? _GEN_515 : _GEN_2358; 
  wire [4:0] _GEN_2441 = integer_inst_r_io_d ? _GEN_516 : _GEN_2359; 
  wire [4:0] _GEN_2442 = integer_inst_r_io_d ? _GEN_517 : _GEN_2360; 
  wire [4:0] _GEN_2443 = integer_inst_r_io_d ? _GEN_518 : _GEN_2361; 
  wire [4:0] _GEN_2444 = integer_inst_r_io_d ? _GEN_519 : _GEN_2362; 
  wire [4:0] _GEN_2445 = integer_inst_r_io_d ? _GEN_520 : _GEN_2363; 
  wire [4:0] _GEN_2446 = integer_inst_r_io_d ? _GEN_521 : _GEN_2364; 
  wire [4:0] _GEN_2447 = integer_inst_r_io_d ? _GEN_522 : _GEN_2365; 
  wire [4:0] _GEN_2448 = integer_inst_r_io_d ? _GEN_523 : _GEN_2366; 
  wire [4:0] _GEN_2449 = integer_inst_r_io_d ? _GEN_524 : _GEN_2367; 
  wire [4:0] _GEN_2450 = integer_inst_r_io_d ? _GEN_525 : _GEN_2368; 
  wire [4:0] _GEN_2451 = integer_inst_r_io_d ? _GEN_526 : _GEN_2369; 
  wire [4:0] _GEN_2452 = integer_inst_r_io_d ? _GEN_527 : _GEN_2370; 
  wire [4:0] _GEN_2453 = integer_inst_r_io_d ? _GEN_528 : _GEN_2371; 
  wire [4:0] _GEN_2454 = integer_inst_r_io_d ? _GEN_529 : _GEN_2372; 
  wire [4:0] _GEN_2455 = integer_inst_r_io_d ? _GEN_530 : _GEN_2373; 
  wire [4:0] _GEN_2456 = integer_inst_r_io_d ? _GEN_531 : _GEN_2374; 
  wire [4:0] _GEN_2457 = integer_inst_r_io_d ? _GEN_532 : _GEN_2375; 
  wire  _GEN_2458 = integer_inst_r_io_d ? _GEN_533 : _GEN_2376; 
  wire  _GEN_2459 = integer_inst_r_io_d ? _GEN_534 : _GEN_2377; 
  wire  _GEN_2460 = integer_inst_r_io_d ? _GEN_535 : _GEN_2378; 
  wire  _GEN_2461 = integer_inst_r_io_d ? _GEN_536 : _GEN_2379; 
  wire  _GEN_2462 = integer_inst_r_io_d ? _GEN_537 : _GEN_2380; 
  wire  _GEN_2463 = integer_inst_r_io_d ? _GEN_538 : _GEN_2381; 
  wire  _GEN_2464 = integer_inst_r_io_d ? _GEN_539 : _GEN_2382; 
  wire  _GEN_2465 = integer_inst_r_io_d ? _GEN_540 : _GEN_2383; 
  wire  _GEN_2466 = integer_inst_r_io_d ? _GEN_541 : _GEN_2384; 
  wire  _GEN_2467 = integer_inst_r_io_d ? _GEN_542 : _GEN_2385; 
  wire  _GEN_2468 = integer_inst_r_io_d ? _GEN_543 : _GEN_2386; 
  wire  _GEN_2469 = integer_inst_r_io_d ? _GEN_544 : _GEN_2387; 
  wire  _GEN_2470 = integer_inst_r_io_d ? _GEN_545 : _GEN_2388; 
  wire  _GEN_2471 = integer_inst_r_io_d ? _GEN_546 : _GEN_2389; 
  wire  _GEN_2472 = integer_inst_r_io_d ? _GEN_547 : _GEN_2390; 
  wire  _GEN_2473 = integer_inst_r_io_d ? _GEN_548 : _GEN_2391; 
  wire  _GEN_2474 = integer_inst_r_io_d ? _GEN_549 : _GEN_2392; 
  wire  _GEN_2475 = integer_inst_r_io_d ? _GEN_550 : _GEN_2393; 
  wire  _GEN_2476 = integer_inst_r_io_d ? _GEN_551 : _GEN_2394; 
  wire  _GEN_2477 = integer_inst_r_io_d ? _GEN_552 : _GEN_2395; 
  wire  _GEN_2478 = integer_inst_r_io_d ? _GEN_553 : _GEN_2396; 
  wire  _GEN_2479 = integer_inst_r_io_d ? _GEN_554 : _GEN_2397; 
  wire  _GEN_2480 = integer_inst_r_io_d ? _GEN_555 : _GEN_2398; 
  wire  _GEN_2481 = integer_inst_r_io_d ? _GEN_556 : _GEN_2399; 
  wire  _GEN_2482 = integer_inst_r_io_d ? _GEN_557 : _GEN_2400; 
  wire  _GEN_2483 = integer_inst_r_io_d ? _GEN_558 : _GEN_2401; 
  wire  _GEN_2484 = integer_inst_r_io_d ? _GEN_559 : _GEN_2402; 
  wire  _GEN_2485 = integer_inst_r_io_d ? _GEN_560 : _GEN_2403; 
  wire  _GEN_2486 = integer_inst_r_io_d ? _GEN_561 : _GEN_2404; 
  wire  _GEN_2487 = integer_inst_r_io_d ? _GEN_562 : _GEN_2405; 
  wire  _GEN_2488 = integer_inst_r_io_d ? _GEN_563 : _GEN_2406; 
  wire  _GEN_2489 = integer_inst_r_io_d ? _GEN_564 : _GEN_2407; 
  wire  _uMulDivOp_io_in_valid_T_1 = uMulDivRS_io_deq_data_qj == 5'h0; 
  wire  _uMulDivOp_io_in_valid_T_2 = ~uMulDivRS__io_empty & _uMulDivOp_io_in_valid_T_1; 
  wire  _uMulDivOp_io_in_valid_T_3 = uMulDivRS_io_deq_data_qk == 5'h0; 
  wire  _uMulDivOp_io_in_valid_T_4 = _uMulDivOp_io_in_valid_T_2 & _uMulDivOp_io_in_valid_T_3; 
  wire  _uMulDivOp_io_in_valid_T_6 = ~uMulDivBusGetData_st_io_q | uCDB_io_muldiv_ready; 
  wire  _rob_addr_match_1_T_2 = uROB_io_queue_data_split_1_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_1 = uROB_io_queue_data_split_1_rob_type == 2'h3 & _rob_addr_match_1_T_2; 
  wire  _rob_addr_match_2_T_2 = uROB_io_queue_data_split_2_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_2 = uROB_io_queue_data_split_2_rob_type == 2'h3 & _rob_addr_match_2_T_2; 
  wire  _rob_addr_match_3_T_2 = uROB_io_queue_data_split_3_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_3 = uROB_io_queue_data_split_3_rob_type == 2'h3 & _rob_addr_match_3_T_2; 
  wire  _rob_addr_match_4_T_2 = uROB_io_queue_data_split_4_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_4 = uROB_io_queue_data_split_4_rob_type == 2'h3 & _rob_addr_match_4_T_2; 
  wire  _rob_addr_match_5_T_2 = uROB_io_queue_data_split_5_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_5 = uROB_io_queue_data_split_5_rob_type == 2'h3 & _rob_addr_match_5_T_2; 
  wire  _rob_addr_match_6_T_2 = uROB_io_queue_data_split_6_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_6 = uROB_io_queue_data_split_6_rob_type == 2'h3 & _rob_addr_match_6_T_2; 
  wire  _rob_addr_match_7_T_2 = uROB_io_queue_data_split_7_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_7 = uROB_io_queue_data_split_7_rob_type == 2'h3 & _rob_addr_match_7_T_2; 
  wire  _rob_addr_match_8_T_2 = uROB_io_queue_data_split_8_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_8 = uROB_io_queue_data_split_8_rob_type == 2'h3 & _rob_addr_match_8_T_2; 
  wire  _rob_addr_match_9_T_2 = uROB_io_queue_data_split_9_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_9 = uROB_io_queue_data_split_9_rob_type == 2'h3 & _rob_addr_match_9_T_2; 
  wire  _rob_addr_match_10_T_2 = uROB_io_queue_data_split_10_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_10 = uROB_io_queue_data_split_10_rob_type == 2'h3 & _rob_addr_match_10_T_2; 
  wire  _rob_addr_match_11_T_2 = uROB_io_queue_data_split_11_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_11 = uROB_io_queue_data_split_11_rob_type == 2'h3 & _rob_addr_match_11_T_2; 
  wire  _rob_addr_match_12_T_2 = uROB_io_queue_data_split_12_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_12 = uROB_io_queue_data_split_12_rob_type == 2'h3 & _rob_addr_match_12_T_2; 
  wire  _rob_addr_match_13_T_2 = uROB_io_queue_data_split_13_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_13 = uROB_io_queue_data_split_13_rob_type == 2'h3 & _rob_addr_match_13_T_2; 
  wire  _rob_addr_match_14_T_2 = uROB_io_queue_data_split_14_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_14 = uROB_io_queue_data_split_14_rob_type == 2'h3 & _rob_addr_match_14_T_2; 
  wire  _rob_addr_match_15_T_2 = uROB_io_queue_data_split_15_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_15 = uROB_io_queue_data_split_15_rob_type == 2'h3 & _rob_addr_match_15_T_2; 
  wire  _rob_addr_match_16_T_2 = uROB_io_queue_data_split_16_rob_dest == issue_mem_addr; 
  wire  rob_addr_match_16 = uROB_io_queue_data_split_16_rob_type == 2'h3 & _rob_addr_match_16_T_2; 
  wire [7:0] addr_match_lo = {rob_addr_match_7,rob_addr_match_6,rob_addr_match_5,rob_addr_match_4,rob_addr_match_3,
    rob_addr_match_2,rob_addr_match_1,1'h0}; 
  wire [16:0] _addr_match_T = {rob_addr_match_16,rob_addr_match_15,rob_addr_match_14,rob_addr_match_13,rob_addr_match_12
    ,rob_addr_match_11,rob_addr_match_10,rob_addr_match_9,rob_addr_match_8,addr_match_lo}; 
  wire  addr_match = |_addr_match_T; 
  wire  uLoadstoreRS_deq_data_op_load = uLoadStoreRS_io_deq_data_op[18]; 
  wire  _datamem_if_ld_valid_T_4 = ~uLoadBusGetData_st_io_q | uCDB_io_mem_ready; 
  wire  _T_634 = ~uROB_io_deq_data_rob_value[0] & uROB__io_deq; 
  wire  _T_637 = uROB_io_deq_data_rob_type == 2'h3; 
  wire [31:0] _GEN_2978 = uROB_io_deq_data_rob_type == 2'h2 ? uROB_io_deq_data_rob_dest : re_jump_addr_r_io_q; 
  wire  _GEN_2979 = uROB_io_deq_data_rob_type == 2'h2 & _T_634; 
  wire  _GEN_2980 = uROB_io_deq_data_rob_type == 2'h2 ? 1'h0 : _T_637; 
  wire  _T_643 = uROB_io_deq_data_rob_dest[5:0] == 6'h1; 
  wire  _T_644 = _T_62 & _T_643; 
  wire  _T_650 = uROB_io_deq_data_rob_dest[5:0] == 6'h2; 
  wire  _T_651 = _T_62 & _T_650; 
  wire  _T_657 = uROB_io_deq_data_rob_dest[5:0] == 6'h3; 
  wire  _T_658 = _T_62 & _T_657; 
  wire  _T_664 = uROB_io_deq_data_rob_dest[5:0] == 6'h4; 
  wire  _T_665 = _T_62 & _T_664; 
  wire  _T_671 = uROB_io_deq_data_rob_dest[5:0] == 6'h5; 
  wire  _T_672 = _T_62 & _T_671; 
  wire  _T_678 = uROB_io_deq_data_rob_dest[5:0] == 6'h6; 
  wire  _T_679 = _T_62 & _T_678; 
  wire  _T_685 = uROB_io_deq_data_rob_dest[5:0] == 6'h7; 
  wire  _T_686 = _T_62 & _T_685; 
  wire  _T_692 = uROB_io_deq_data_rob_dest[5:0] == 6'h8; 
  wire  _T_693 = _T_62 & _T_692; 
  wire  _T_699 = uROB_io_deq_data_rob_dest[5:0] == 6'h9; 
  wire  _T_700 = _T_62 & _T_699; 
  wire  _T_706 = uROB_io_deq_data_rob_dest[5:0] == 6'ha; 
  wire  _T_707 = _T_62 & _T_706; 
  wire  _T_713 = uROB_io_deq_data_rob_dest[5:0] == 6'hb; 
  wire  _T_714 = _T_62 & _T_713; 
  wire  _T_720 = uROB_io_deq_data_rob_dest[5:0] == 6'hc; 
  wire  _T_721 = _T_62 & _T_720; 
  wire  _T_727 = uROB_io_deq_data_rob_dest[5:0] == 6'hd; 
  wire  _T_728 = _T_62 & _T_727; 
  wire  _T_734 = uROB_io_deq_data_rob_dest[5:0] == 6'he; 
  wire  _T_735 = _T_62 & _T_734; 
  wire  _T_741 = uROB_io_deq_data_rob_dest[5:0] == 6'hf; 
  wire  _T_742 = _T_62 & _T_741; 
  wire  _T_748 = uROB_io_deq_data_rob_dest[5:0] == 6'h10; 
  wire  _T_749 = _T_62 & _T_748; 
  wire  _T_755 = uROB_io_deq_data_rob_dest[5:0] == 6'h11; 
  wire  _T_756 = _T_62 & _T_755; 
  wire  _T_762 = uROB_io_deq_data_rob_dest[5:0] == 6'h12; 
  wire  _T_763 = _T_62 & _T_762; 
  wire  _T_769 = uROB_io_deq_data_rob_dest[5:0] == 6'h13; 
  wire  _T_770 = _T_62 & _T_769; 
  wire  _T_776 = uROB_io_deq_data_rob_dest[5:0] == 6'h14; 
  wire  _T_777 = _T_62 & _T_776; 
  wire  _T_783 = uROB_io_deq_data_rob_dest[5:0] == 6'h15; 
  wire  _T_784 = _T_62 & _T_783; 
  wire  _T_790 = uROB_io_deq_data_rob_dest[5:0] == 6'h16; 
  wire  _T_791 = _T_62 & _T_790; 
  wire  _T_797 = uROB_io_deq_data_rob_dest[5:0] == 6'h17; 
  wire  _T_798 = _T_62 & _T_797; 
  wire  _T_804 = uROB_io_deq_data_rob_dest[5:0] == 6'h18; 
  wire  _T_805 = _T_62 & _T_804; 
  wire  _T_811 = uROB_io_deq_data_rob_dest[5:0] == 6'h19; 
  wire  _T_812 = _T_62 & _T_811; 
  wire  _T_818 = uROB_io_deq_data_rob_dest[5:0] == 6'h1a; 
  wire  _T_819 = _T_62 & _T_818; 
  wire  _T_825 = uROB_io_deq_data_rob_dest[5:0] == 6'h1b; 
  wire  _T_826 = _T_62 & _T_825; 
  wire  _T_832 = uROB_io_deq_data_rob_dest[5:0] == 6'h1c; 
  wire  _T_833 = _T_62 & _T_832; 
  wire  _T_839 = uROB_io_deq_data_rob_dest[5:0] == 6'h1d; 
  wire  _T_840 = _T_62 & _T_839; 
  wire  _T_846 = uROB_io_deq_data_rob_dest[5:0] == 6'h1e; 
  wire  _T_847 = _T_62 & _T_846; 
  wire  _T_853 = uROB_io_deq_data_rob_dest[5:0] == 6'h1f; 
  wire  _T_854 = _T_62 & _T_853; 
  integer_RS uIntergerRS_ ( 
    .clock(uIntergerRS__clock),
    .reset(uIntergerRS__reset),
    .io_clear(uIntergerRS__io_clear),
    .io_enq(uIntergerRS__io_enq),
    .io_enq_data(uIntergerRS__io_enq_data),
    .io_deq(uIntergerRS__io_deq),
    .io_deq_cond(uIntergerRS__io_deq_cond),
    .io_deq_data(uIntergerRS__io_deq_data),
    .io_empty(uIntergerRS__io_empty),
    .io_full(uIntergerRS__io_full),
    .io_queue_data(uIntergerRS__io_queue_data),
    .io_update_entry(uIntergerRS__io_update_entry),
    .io_update_entry_data(uIntergerRS__io_update_entry_data)
  );
  FIFO uMulDivRS_ ( 
    .clock(uMulDivRS__clock),
    .reset(uMulDivRS__reset),
    .io_clear(uMulDivRS__io_clear),
    .io_enq(uMulDivRS__io_enq),
    .io_enq_data(uMulDivRS__io_enq_data),
    .io_enq_idx(uMulDivRS__io_enq_idx),
    .io_deq(uMulDivRS__io_deq),
    .io_deq_data(uMulDivRS__io_deq_data),
    .io_deq_idx(uMulDivRS__io_deq_idx),
    .io_empty(uMulDivRS__io_empty),
    .io_full(uMulDivRS__io_full),
    .io_queue_data(uMulDivRS__io_queue_data),
    .io_update_entry(uMulDivRS__io_update_entry),
    .io_update_entry_data(uMulDivRS__io_update_entry_data)
  );
  FIFO uLoadStoreRS_ ( 
    .clock(uLoadStoreRS__clock),
    .reset(uLoadStoreRS__reset),
    .io_clear(uLoadStoreRS__io_clear),
    .io_enq(uLoadStoreRS__io_enq),
    .io_enq_data(uLoadStoreRS__io_enq_data),
    .io_enq_idx(uLoadStoreRS__io_enq_idx),
    .io_deq(uLoadStoreRS__io_deq),
    .io_deq_data(uLoadStoreRS__io_deq_data),
    .io_deq_idx(uLoadStoreRS__io_deq_idx),
    .io_empty(uLoadStoreRS__io_empty),
    .io_full(uLoadStoreRS__io_full),
    .io_queue_data(uLoadStoreRS__io_queue_data),
    .io_update_entry(uLoadStoreRS__io_update_entry),
    .io_update_entry_data(uLoadStoreRS__io_update_entry_data)
  );
  FIFO_ROB uROB_ ( 
    .clock(uROB__clock),
    .reset(uROB__reset),
    .io_clear(uROB__io_clear),
    .io_enq(uROB__io_enq),
    .io_enq_data(uROB__io_enq_data),
    .io_deq(uROB__io_deq),
    .io_deq_data(uROB__io_deq_data),
    .io_empty(uROB__io_empty),
    .io_full(uROB__io_full),
    .io_enq_idx(uROB__io_enq_idx),
    .io_deq_idx(uROB__io_deq_idx),
    .io_queue_data(uROB__io_queue_data),
    .io_update_entry(uROB__io_update_entry),
    .io_update_entry_data(uROB__io_update_entry_data)
  );
  CDB uCDB ( 
    .clock(uCDB_clock),
    .reset(uCDB_reset),
    .io_clear(uCDB_io_clear),
    .io_int_valid(uCDB_io_int_valid),
    .io_int_ready(uCDB_io_int_ready),
    .io_int_result(uCDB_io_int_result),
    .io_int_dest(uCDB_io_int_dest),
    .io_muldiv_valid(uCDB_io_muldiv_valid),
    .io_muldiv_ready(uCDB_io_muldiv_ready),
    .io_muldiv_result(uCDB_io_muldiv_result),
    .io_muldiv_dest(uCDB_io_muldiv_dest),
    .io_mem_valid(uCDB_io_mem_valid),
    .io_mem_ready(uCDB_io_mem_ready),
    .io_mem_result(uCDB_io_mem_result),
    .io_mem_dest(uCDB_io_mem_dest),
    .io_cdb_valid(uCDB_io_cdb_valid),
    .io_cdb_result(uCDB_io_cdb_result),
    .io_cdb_dest(uCDB_io_cdb_dest)
  );
  IntOp uIntOp ( 
    .clock(uIntOp_clock),
    .reset(uIntOp_reset),
    .io_clear(uIntOp_io_clear),
    .io_in_valid(uIntOp_io_in_valid),
    .io_in_in1(uIntOp_io_in_in1),
    .io_in_in2(uIntOp_io_in_in2),
    .io_in_op_store(uIntOp_io_in_op_store),
    .io_in_op_load(uIntOp_io_in_op_load),
    .io_in_op_muldivb_s(uIntOp_io_in_op_muldivb_s),
    .io_in_op_muldiva_s(uIntOp_io_in_op_muldiva_s),
    .io_in_op_div(uIntOp_io_in_op_div),
    .io_in_op_mul(uIntOp_io_in_op_mul),
    .io_in_op_equal(uIntOp_io_in_op_equal),
    .io_in_op_large(uIntOp_io_in_op_large),
    .io_in_op_less(uIntOp_io_in_op_less),
    .io_in_op_jr(uIntOp_io_in_op_jr),
    .io_in_op_br(uIntOp_io_in_op_br),
    .io_in_op_sra(uIntOp_io_in_op_sra),
    .io_in_op_srl(uIntOp_io_in_op_srl),
    .io_in_op_sll(uIntOp_io_in_op_sll),
    .io_in_op_sub(uIntOp_io_in_op_sub),
    .io_in_op_add(uIntOp_io_in_op_add),
    .io_in_op_set(uIntOp_io_in_op_set),
    .io_in_op_xor(uIntOp_io_in_op_xor),
    .io_in_op_or(uIntOp_io_in_op_or),
    .io_in_op_and(uIntOp_io_in_op_and),
    .io_in_dest(uIntOp_io_in_dest),
    .io_out_valid(uIntOp_io_out_valid),
    .io_out_result(uIntOp_io_out_result),
    .io_out_dest(uIntOp_io_out_dest)
  );
  MulDivOp uMulDivOp ( 
    .clock(uMulDivOp_clock),
    .reset(uMulDivOp_reset),
    .io_clear(uMulDivOp_io_clear),
    .io_in_valid(uMulDivOp_io_in_valid),
    .io_in_in1(uMulDivOp_io_in_in1),
    .io_in_in2(uMulDivOp_io_in_in2),
    .io_in_op_muldivb_s(uMulDivOp_io_in_op_muldivb_s),
    .io_in_op_muldiva_s(uMulDivOp_io_in_op_muldiva_s),
    .io_in_op_mul(uMulDivOp_io_in_op_mul),
    .io_in_dest(uMulDivOp_io_in_dest),
    .io_out_valid(uMulDivOp_io_out_valid),
    .io_out_result(uMulDivOp_io_out_result),
    .io_out_dest(uMulDivOp_io_out_dest)
  );
  prim_ff_cl_39 uRegFile_0 ( 
    .clock(uRegFile_0_clock),
    .reset(uRegFile_0_reset),
    .io_q(uRegFile_0_io_q),
    .io_d(uRegFile_0_io_d),
    .io_clear(uRegFile_0_io_clear)
  );
  prim_ff_cl_39 uRegFile_1 ( 
    .clock(uRegFile_1_clock),
    .reset(uRegFile_1_reset),
    .io_q(uRegFile_1_io_q),
    .io_d(uRegFile_1_io_d),
    .io_clear(uRegFile_1_io_clear)
  );
  prim_ff_cl_39 uRegFile_2 ( 
    .clock(uRegFile_2_clock),
    .reset(uRegFile_2_reset),
    .io_q(uRegFile_2_io_q),
    .io_d(uRegFile_2_io_d),
    .io_clear(uRegFile_2_io_clear)
  );
  prim_ff_cl_39 uRegFile_3 ( 
    .clock(uRegFile_3_clock),
    .reset(uRegFile_3_reset),
    .io_q(uRegFile_3_io_q),
    .io_d(uRegFile_3_io_d),
    .io_clear(uRegFile_3_io_clear)
  );
  prim_ff_cl_39 uRegFile_4 ( 
    .clock(uRegFile_4_clock),
    .reset(uRegFile_4_reset),
    .io_q(uRegFile_4_io_q),
    .io_d(uRegFile_4_io_d),
    .io_clear(uRegFile_4_io_clear)
  );
  prim_ff_cl_39 uRegFile_5 ( 
    .clock(uRegFile_5_clock),
    .reset(uRegFile_5_reset),
    .io_q(uRegFile_5_io_q),
    .io_d(uRegFile_5_io_d),
    .io_clear(uRegFile_5_io_clear)
  );
  prim_ff_cl_39 uRegFile_6 ( 
    .clock(uRegFile_6_clock),
    .reset(uRegFile_6_reset),
    .io_q(uRegFile_6_io_q),
    .io_d(uRegFile_6_io_d),
    .io_clear(uRegFile_6_io_clear)
  );
  prim_ff_cl_39 uRegFile_7 ( 
    .clock(uRegFile_7_clock),
    .reset(uRegFile_7_reset),
    .io_q(uRegFile_7_io_q),
    .io_d(uRegFile_7_io_d),
    .io_clear(uRegFile_7_io_clear)
  );
  prim_ff_cl_39 uRegFile_8 ( 
    .clock(uRegFile_8_clock),
    .reset(uRegFile_8_reset),
    .io_q(uRegFile_8_io_q),
    .io_d(uRegFile_8_io_d),
    .io_clear(uRegFile_8_io_clear)
  );
  prim_ff_cl_39 uRegFile_9 ( 
    .clock(uRegFile_9_clock),
    .reset(uRegFile_9_reset),
    .io_q(uRegFile_9_io_q),
    .io_d(uRegFile_9_io_d),
    .io_clear(uRegFile_9_io_clear)
  );
  prim_ff_cl_39 uRegFile_10 ( 
    .clock(uRegFile_10_clock),
    .reset(uRegFile_10_reset),
    .io_q(uRegFile_10_io_q),
    .io_d(uRegFile_10_io_d),
    .io_clear(uRegFile_10_io_clear)
  );
  prim_ff_cl_39 uRegFile_11 ( 
    .clock(uRegFile_11_clock),
    .reset(uRegFile_11_reset),
    .io_q(uRegFile_11_io_q),
    .io_d(uRegFile_11_io_d),
    .io_clear(uRegFile_11_io_clear)
  );
  prim_ff_cl_39 uRegFile_12 ( 
    .clock(uRegFile_12_clock),
    .reset(uRegFile_12_reset),
    .io_q(uRegFile_12_io_q),
    .io_d(uRegFile_12_io_d),
    .io_clear(uRegFile_12_io_clear)
  );
  prim_ff_cl_39 uRegFile_13 ( 
    .clock(uRegFile_13_clock),
    .reset(uRegFile_13_reset),
    .io_q(uRegFile_13_io_q),
    .io_d(uRegFile_13_io_d),
    .io_clear(uRegFile_13_io_clear)
  );
  prim_ff_cl_39 uRegFile_14 ( 
    .clock(uRegFile_14_clock),
    .reset(uRegFile_14_reset),
    .io_q(uRegFile_14_io_q),
    .io_d(uRegFile_14_io_d),
    .io_clear(uRegFile_14_io_clear)
  );
  prim_ff_cl_39 uRegFile_15 ( 
    .clock(uRegFile_15_clock),
    .reset(uRegFile_15_reset),
    .io_q(uRegFile_15_io_q),
    .io_d(uRegFile_15_io_d),
    .io_clear(uRegFile_15_io_clear)
  );
  prim_ff_cl_39 uRegFile_16 ( 
    .clock(uRegFile_16_clock),
    .reset(uRegFile_16_reset),
    .io_q(uRegFile_16_io_q),
    .io_d(uRegFile_16_io_d),
    .io_clear(uRegFile_16_io_clear)
  );
  prim_ff_cl_39 uRegFile_17 ( 
    .clock(uRegFile_17_clock),
    .reset(uRegFile_17_reset),
    .io_q(uRegFile_17_io_q),
    .io_d(uRegFile_17_io_d),
    .io_clear(uRegFile_17_io_clear)
  );
  prim_ff_cl_39 uRegFile_18 ( 
    .clock(uRegFile_18_clock),
    .reset(uRegFile_18_reset),
    .io_q(uRegFile_18_io_q),
    .io_d(uRegFile_18_io_d),
    .io_clear(uRegFile_18_io_clear)
  );
  prim_ff_cl_39 uRegFile_19 ( 
    .clock(uRegFile_19_clock),
    .reset(uRegFile_19_reset),
    .io_q(uRegFile_19_io_q),
    .io_d(uRegFile_19_io_d),
    .io_clear(uRegFile_19_io_clear)
  );
  prim_ff_cl_39 uRegFile_20 ( 
    .clock(uRegFile_20_clock),
    .reset(uRegFile_20_reset),
    .io_q(uRegFile_20_io_q),
    .io_d(uRegFile_20_io_d),
    .io_clear(uRegFile_20_io_clear)
  );
  prim_ff_cl_39 uRegFile_21 ( 
    .clock(uRegFile_21_clock),
    .reset(uRegFile_21_reset),
    .io_q(uRegFile_21_io_q),
    .io_d(uRegFile_21_io_d),
    .io_clear(uRegFile_21_io_clear)
  );
  prim_ff_cl_39 uRegFile_22 ( 
    .clock(uRegFile_22_clock),
    .reset(uRegFile_22_reset),
    .io_q(uRegFile_22_io_q),
    .io_d(uRegFile_22_io_d),
    .io_clear(uRegFile_22_io_clear)
  );
  prim_ff_cl_39 uRegFile_23 ( 
    .clock(uRegFile_23_clock),
    .reset(uRegFile_23_reset),
    .io_q(uRegFile_23_io_q),
    .io_d(uRegFile_23_io_d),
    .io_clear(uRegFile_23_io_clear)
  );
  prim_ff_cl_39 uRegFile_24 ( 
    .clock(uRegFile_24_clock),
    .reset(uRegFile_24_reset),
    .io_q(uRegFile_24_io_q),
    .io_d(uRegFile_24_io_d),
    .io_clear(uRegFile_24_io_clear)
  );
  prim_ff_cl_39 uRegFile_25 ( 
    .clock(uRegFile_25_clock),
    .reset(uRegFile_25_reset),
    .io_q(uRegFile_25_io_q),
    .io_d(uRegFile_25_io_d),
    .io_clear(uRegFile_25_io_clear)
  );
  prim_ff_cl_39 uRegFile_26 ( 
    .clock(uRegFile_26_clock),
    .reset(uRegFile_26_reset),
    .io_q(uRegFile_26_io_q),
    .io_d(uRegFile_26_io_d),
    .io_clear(uRegFile_26_io_clear)
  );
  prim_ff_cl_39 uRegFile_27 ( 
    .clock(uRegFile_27_clock),
    .reset(uRegFile_27_reset),
    .io_q(uRegFile_27_io_q),
    .io_d(uRegFile_27_io_d),
    .io_clear(uRegFile_27_io_clear)
  );
  prim_ff_cl_39 uRegFile_28 ( 
    .clock(uRegFile_28_clock),
    .reset(uRegFile_28_reset),
    .io_q(uRegFile_28_io_q),
    .io_d(uRegFile_28_io_d),
    .io_clear(uRegFile_28_io_clear)
  );
  prim_ff_cl_39 uRegFile_29 ( 
    .clock(uRegFile_29_clock),
    .reset(uRegFile_29_reset),
    .io_q(uRegFile_29_io_q),
    .io_d(uRegFile_29_io_d),
    .io_clear(uRegFile_29_io_clear)
  );
  prim_ff_cl_39 uRegFile_30 ( 
    .clock(uRegFile_30_clock),
    .reset(uRegFile_30_reset),
    .io_q(uRegFile_30_io_q),
    .io_d(uRegFile_30_io_d),
    .io_clear(uRegFile_30_io_clear)
  );
  prim_ff_cl_39 uRegFile_31 ( 
    .clock(uRegFile_31_clock),
    .reset(uRegFile_31_reset),
    .io_q(uRegFile_31_io_q),
    .io_d(uRegFile_31_io_d),
    .io_clear(uRegFile_31_io_clear)
  );
  prim_ff_cl_71 uRegState_0 ( 
    .clock(uRegState_0_clock),
    .reset(uRegState_0_reset),
    .io_q_busy(uRegState_0_io_q_busy),
    .io_q_reorder(uRegState_0_io_q_reorder),
    .io_d_busy(uRegState_0_io_d_busy),
    .io_d_reorder(uRegState_0_io_d_reorder),
    .io_clear(uRegState_0_io_clear)
  );
  prim_ff_cl_71 uRegState_1 ( 
    .clock(uRegState_1_clock),
    .reset(uRegState_1_reset),
    .io_q_busy(uRegState_1_io_q_busy),
    .io_q_reorder(uRegState_1_io_q_reorder),
    .io_d_busy(uRegState_1_io_d_busy),
    .io_d_reorder(uRegState_1_io_d_reorder),
    .io_clear(uRegState_1_io_clear)
  );
  prim_ff_cl_71 uRegState_2 ( 
    .clock(uRegState_2_clock),
    .reset(uRegState_2_reset),
    .io_q_busy(uRegState_2_io_q_busy),
    .io_q_reorder(uRegState_2_io_q_reorder),
    .io_d_busy(uRegState_2_io_d_busy),
    .io_d_reorder(uRegState_2_io_d_reorder),
    .io_clear(uRegState_2_io_clear)
  );
  prim_ff_cl_71 uRegState_3 ( 
    .clock(uRegState_3_clock),
    .reset(uRegState_3_reset),
    .io_q_busy(uRegState_3_io_q_busy),
    .io_q_reorder(uRegState_3_io_q_reorder),
    .io_d_busy(uRegState_3_io_d_busy),
    .io_d_reorder(uRegState_3_io_d_reorder),
    .io_clear(uRegState_3_io_clear)
  );
  prim_ff_cl_71 uRegState_4 ( 
    .clock(uRegState_4_clock),
    .reset(uRegState_4_reset),
    .io_q_busy(uRegState_4_io_q_busy),
    .io_q_reorder(uRegState_4_io_q_reorder),
    .io_d_busy(uRegState_4_io_d_busy),
    .io_d_reorder(uRegState_4_io_d_reorder),
    .io_clear(uRegState_4_io_clear)
  );
  prim_ff_cl_71 uRegState_5 ( 
    .clock(uRegState_5_clock),
    .reset(uRegState_5_reset),
    .io_q_busy(uRegState_5_io_q_busy),
    .io_q_reorder(uRegState_5_io_q_reorder),
    .io_d_busy(uRegState_5_io_d_busy),
    .io_d_reorder(uRegState_5_io_d_reorder),
    .io_clear(uRegState_5_io_clear)
  );
  prim_ff_cl_71 uRegState_6 ( 
    .clock(uRegState_6_clock),
    .reset(uRegState_6_reset),
    .io_q_busy(uRegState_6_io_q_busy),
    .io_q_reorder(uRegState_6_io_q_reorder),
    .io_d_busy(uRegState_6_io_d_busy),
    .io_d_reorder(uRegState_6_io_d_reorder),
    .io_clear(uRegState_6_io_clear)
  );
  prim_ff_cl_71 uRegState_7 ( 
    .clock(uRegState_7_clock),
    .reset(uRegState_7_reset),
    .io_q_busy(uRegState_7_io_q_busy),
    .io_q_reorder(uRegState_7_io_q_reorder),
    .io_d_busy(uRegState_7_io_d_busy),
    .io_d_reorder(uRegState_7_io_d_reorder),
    .io_clear(uRegState_7_io_clear)
  );
  prim_ff_cl_71 uRegState_8 ( 
    .clock(uRegState_8_clock),
    .reset(uRegState_8_reset),
    .io_q_busy(uRegState_8_io_q_busy),
    .io_q_reorder(uRegState_8_io_q_reorder),
    .io_d_busy(uRegState_8_io_d_busy),
    .io_d_reorder(uRegState_8_io_d_reorder),
    .io_clear(uRegState_8_io_clear)
  );
  prim_ff_cl_71 uRegState_9 ( 
    .clock(uRegState_9_clock),
    .reset(uRegState_9_reset),
    .io_q_busy(uRegState_9_io_q_busy),
    .io_q_reorder(uRegState_9_io_q_reorder),
    .io_d_busy(uRegState_9_io_d_busy),
    .io_d_reorder(uRegState_9_io_d_reorder),
    .io_clear(uRegState_9_io_clear)
  );
  prim_ff_cl_71 uRegState_10 ( 
    .clock(uRegState_10_clock),
    .reset(uRegState_10_reset),
    .io_q_busy(uRegState_10_io_q_busy),
    .io_q_reorder(uRegState_10_io_q_reorder),
    .io_d_busy(uRegState_10_io_d_busy),
    .io_d_reorder(uRegState_10_io_d_reorder),
    .io_clear(uRegState_10_io_clear)
  );
  prim_ff_cl_71 uRegState_11 ( 
    .clock(uRegState_11_clock),
    .reset(uRegState_11_reset),
    .io_q_busy(uRegState_11_io_q_busy),
    .io_q_reorder(uRegState_11_io_q_reorder),
    .io_d_busy(uRegState_11_io_d_busy),
    .io_d_reorder(uRegState_11_io_d_reorder),
    .io_clear(uRegState_11_io_clear)
  );
  prim_ff_cl_71 uRegState_12 ( 
    .clock(uRegState_12_clock),
    .reset(uRegState_12_reset),
    .io_q_busy(uRegState_12_io_q_busy),
    .io_q_reorder(uRegState_12_io_q_reorder),
    .io_d_busy(uRegState_12_io_d_busy),
    .io_d_reorder(uRegState_12_io_d_reorder),
    .io_clear(uRegState_12_io_clear)
  );
  prim_ff_cl_71 uRegState_13 ( 
    .clock(uRegState_13_clock),
    .reset(uRegState_13_reset),
    .io_q_busy(uRegState_13_io_q_busy),
    .io_q_reorder(uRegState_13_io_q_reorder),
    .io_d_busy(uRegState_13_io_d_busy),
    .io_d_reorder(uRegState_13_io_d_reorder),
    .io_clear(uRegState_13_io_clear)
  );
  prim_ff_cl_71 uRegState_14 ( 
    .clock(uRegState_14_clock),
    .reset(uRegState_14_reset),
    .io_q_busy(uRegState_14_io_q_busy),
    .io_q_reorder(uRegState_14_io_q_reorder),
    .io_d_busy(uRegState_14_io_d_busy),
    .io_d_reorder(uRegState_14_io_d_reorder),
    .io_clear(uRegState_14_io_clear)
  );
  prim_ff_cl_71 uRegState_15 ( 
    .clock(uRegState_15_clock),
    .reset(uRegState_15_reset),
    .io_q_busy(uRegState_15_io_q_busy),
    .io_q_reorder(uRegState_15_io_q_reorder),
    .io_d_busy(uRegState_15_io_d_busy),
    .io_d_reorder(uRegState_15_io_d_reorder),
    .io_clear(uRegState_15_io_clear)
  );
  prim_ff_cl_71 uRegState_16 ( 
    .clock(uRegState_16_clock),
    .reset(uRegState_16_reset),
    .io_q_busy(uRegState_16_io_q_busy),
    .io_q_reorder(uRegState_16_io_q_reorder),
    .io_d_busy(uRegState_16_io_d_busy),
    .io_d_reorder(uRegState_16_io_d_reorder),
    .io_clear(uRegState_16_io_clear)
  );
  prim_ff_cl_71 uRegState_17 ( 
    .clock(uRegState_17_clock),
    .reset(uRegState_17_reset),
    .io_q_busy(uRegState_17_io_q_busy),
    .io_q_reorder(uRegState_17_io_q_reorder),
    .io_d_busy(uRegState_17_io_d_busy),
    .io_d_reorder(uRegState_17_io_d_reorder),
    .io_clear(uRegState_17_io_clear)
  );
  prim_ff_cl_71 uRegState_18 ( 
    .clock(uRegState_18_clock),
    .reset(uRegState_18_reset),
    .io_q_busy(uRegState_18_io_q_busy),
    .io_q_reorder(uRegState_18_io_q_reorder),
    .io_d_busy(uRegState_18_io_d_busy),
    .io_d_reorder(uRegState_18_io_d_reorder),
    .io_clear(uRegState_18_io_clear)
  );
  prim_ff_cl_71 uRegState_19 ( 
    .clock(uRegState_19_clock),
    .reset(uRegState_19_reset),
    .io_q_busy(uRegState_19_io_q_busy),
    .io_q_reorder(uRegState_19_io_q_reorder),
    .io_d_busy(uRegState_19_io_d_busy),
    .io_d_reorder(uRegState_19_io_d_reorder),
    .io_clear(uRegState_19_io_clear)
  );
  prim_ff_cl_71 uRegState_20 ( 
    .clock(uRegState_20_clock),
    .reset(uRegState_20_reset),
    .io_q_busy(uRegState_20_io_q_busy),
    .io_q_reorder(uRegState_20_io_q_reorder),
    .io_d_busy(uRegState_20_io_d_busy),
    .io_d_reorder(uRegState_20_io_d_reorder),
    .io_clear(uRegState_20_io_clear)
  );
  prim_ff_cl_71 uRegState_21 ( 
    .clock(uRegState_21_clock),
    .reset(uRegState_21_reset),
    .io_q_busy(uRegState_21_io_q_busy),
    .io_q_reorder(uRegState_21_io_q_reorder),
    .io_d_busy(uRegState_21_io_d_busy),
    .io_d_reorder(uRegState_21_io_d_reorder),
    .io_clear(uRegState_21_io_clear)
  );
  prim_ff_cl_71 uRegState_22 ( 
    .clock(uRegState_22_clock),
    .reset(uRegState_22_reset),
    .io_q_busy(uRegState_22_io_q_busy),
    .io_q_reorder(uRegState_22_io_q_reorder),
    .io_d_busy(uRegState_22_io_d_busy),
    .io_d_reorder(uRegState_22_io_d_reorder),
    .io_clear(uRegState_22_io_clear)
  );
  prim_ff_cl_71 uRegState_23 ( 
    .clock(uRegState_23_clock),
    .reset(uRegState_23_reset),
    .io_q_busy(uRegState_23_io_q_busy),
    .io_q_reorder(uRegState_23_io_q_reorder),
    .io_d_busy(uRegState_23_io_d_busy),
    .io_d_reorder(uRegState_23_io_d_reorder),
    .io_clear(uRegState_23_io_clear)
  );
  prim_ff_cl_71 uRegState_24 ( 
    .clock(uRegState_24_clock),
    .reset(uRegState_24_reset),
    .io_q_busy(uRegState_24_io_q_busy),
    .io_q_reorder(uRegState_24_io_q_reorder),
    .io_d_busy(uRegState_24_io_d_busy),
    .io_d_reorder(uRegState_24_io_d_reorder),
    .io_clear(uRegState_24_io_clear)
  );
  prim_ff_cl_71 uRegState_25 ( 
    .clock(uRegState_25_clock),
    .reset(uRegState_25_reset),
    .io_q_busy(uRegState_25_io_q_busy),
    .io_q_reorder(uRegState_25_io_q_reorder),
    .io_d_busy(uRegState_25_io_d_busy),
    .io_d_reorder(uRegState_25_io_d_reorder),
    .io_clear(uRegState_25_io_clear)
  );
  prim_ff_cl_71 uRegState_26 ( 
    .clock(uRegState_26_clock),
    .reset(uRegState_26_reset),
    .io_q_busy(uRegState_26_io_q_busy),
    .io_q_reorder(uRegState_26_io_q_reorder),
    .io_d_busy(uRegState_26_io_d_busy),
    .io_d_reorder(uRegState_26_io_d_reorder),
    .io_clear(uRegState_26_io_clear)
  );
  prim_ff_cl_71 uRegState_27 ( 
    .clock(uRegState_27_clock),
    .reset(uRegState_27_reset),
    .io_q_busy(uRegState_27_io_q_busy),
    .io_q_reorder(uRegState_27_io_q_reorder),
    .io_d_busy(uRegState_27_io_d_busy),
    .io_d_reorder(uRegState_27_io_d_reorder),
    .io_clear(uRegState_27_io_clear)
  );
  prim_ff_cl_71 uRegState_28 ( 
    .clock(uRegState_28_clock),
    .reset(uRegState_28_reset),
    .io_q_busy(uRegState_28_io_q_busy),
    .io_q_reorder(uRegState_28_io_q_reorder),
    .io_d_busy(uRegState_28_io_d_busy),
    .io_d_reorder(uRegState_28_io_d_reorder),
    .io_clear(uRegState_28_io_clear)
  );
  prim_ff_cl_71 uRegState_29 ( 
    .clock(uRegState_29_clock),
    .reset(uRegState_29_reset),
    .io_q_busy(uRegState_29_io_q_busy),
    .io_q_reorder(uRegState_29_io_q_reorder),
    .io_d_busy(uRegState_29_io_d_busy),
    .io_d_reorder(uRegState_29_io_d_reorder),
    .io_clear(uRegState_29_io_clear)
  );
  prim_ff_cl_71 uRegState_30 ( 
    .clock(uRegState_30_clock),
    .reset(uRegState_30_reset),
    .io_q_busy(uRegState_30_io_q_busy),
    .io_q_reorder(uRegState_30_io_q_reorder),
    .io_d_busy(uRegState_30_io_d_busy),
    .io_d_reorder(uRegState_30_io_d_reorder),
    .io_clear(uRegState_30_io_clear)
  );
  prim_ff_cl_71 uRegState_31 ( 
    .clock(uRegState_31_clock),
    .reset(uRegState_31_reset),
    .io_q_busy(uRegState_31_io_q_busy),
    .io_q_reorder(uRegState_31_io_q_reorder),
    .io_d_busy(uRegState_31_io_d_busy),
    .io_d_reorder(uRegState_31_io_d_reorder),
    .io_clear(uRegState_31_io_clear)
  );
  prim_ff_cl_103 integer_inst_r ( 
    .clock(integer_inst_r_clock),
    .reset(integer_inst_r_reset),
    .io_q(integer_inst_r_io_q),
    .io_d(integer_inst_r_io_d),
    .io_clear(integer_inst_r_io_clear)
  );
  prim_ff_cl_103 branch_inst_r ( 
    .clock(branch_inst_r_clock),
    .reset(branch_inst_r_reset),
    .io_q(branch_inst_r_io_q),
    .io_d(branch_inst_r_io_d),
    .io_clear(branch_inst_r_io_clear)
  );
  prim_ff_cl_103 store_inst_r ( 
    .clock(store_inst_r_clock),
    .reset(store_inst_r_reset),
    .io_q(store_inst_r_io_q),
    .io_d(store_inst_r_io_d),
    .io_clear(store_inst_r_io_clear)
  );
  prim_ff_cl_103 load_inst_r ( 
    .clock(load_inst_r_clock),
    .reset(load_inst_r_reset),
    .io_q(load_inst_r_io_q),
    .io_d(load_inst_r_io_d),
    .io_clear(load_inst_r_io_clear)
  );
  prim_ff_cl_103 muldiv_inst_r ( 
    .clock(muldiv_inst_r_clock),
    .reset(muldiv_inst_r_reset),
    .io_q(muldiv_inst_r_io_q),
    .io_d(muldiv_inst_r_io_d),
    .io_clear(muldiv_inst_r_io_clear)
  );
  prim_ff_cl_5 mBranchProc_st ( 
    .clock(mBranchProc_st_clock),
    .reset(mBranchProc_st_reset),
    .io_q(mBranchProc_st_io_q),
    .io_d(mBranchProc_st_io_d),
    .io_clear(mBranchProc_st_io_clear)
  );
  prim_ff_cl_39 re_jump_addr_r ( 
    .clock(re_jump_addr_r_clock),
    .reset(re_jump_addr_r_reset),
    .io_q(re_jump_addr_r_io_q),
    .io_d(re_jump_addr_r_io_d),
    .io_clear(re_jump_addr_r_io_clear)
  );
  prim_ff_cl_103 uIntBusGetData_st ( 
    .clock(uIntBusGetData_st_clock),
    .reset(uIntBusGetData_st_reset),
    .io_q(uIntBusGetData_st_io_q),
    .io_d(uIntBusGetData_st_io_d),
    .io_clear(uIntBusGetData_st_io_clear)
  );
  prim_ff_cl_103 uMulDivBusGetData_st ( 
    .clock(uMulDivBusGetData_st_clock),
    .reset(uMulDivBusGetData_st_reset),
    .io_q(uMulDivBusGetData_st_io_q),
    .io_d(uMulDivBusGetData_st_io_d),
    .io_clear(uMulDivBusGetData_st_io_clear)
  );
  prim_ff_cl_103 uLoadBusGetData_st ( 
    .clock(uLoadBusGetData_st_clock),
    .reset(uLoadBusGetData_st_reset),
    .io_q(uLoadBusGetData_st_io_q),
    .io_d(uLoadBusGetData_st_io_d),
    .io_clear(uLoadBusGetData_st_io_clear)
  );
  assign fetcher_if_stall_fetch = 2'h0 == branchProc_stEnum ? _GEN_12 : _GEN_16; 
  assign fetcher_if_re_jump_en = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign fetcher_if_re_jump_addr = re_jump_addr_r_io_d; 
  assign datamem_if_RS_idx_i = uLoadStoreRS__io_deq_data[111:107]; 
  assign datamem_if_st_valid = uROB_io_deq_data_rob_ready & _GEN_2980; 
  assign datamem_if_st_addr = uROB__io_deq_data[64:33]; 
  assign datamem_if_st_data = uROB__io_deq_data[32:1]; 
  assign datamem_if_ld_valid = ~addr_match & uLoadstoreRS_deq_data_op_load & uLoadStoreRS_out_valid &
    _datamem_if_ld_valid_T_4; 
  assign datamem_if_ld_addr = uLoadStoreRS_io_deq_data_vj + uLoadStoreRS_io_deq_data_a; 
  assign uIntergerRS__clock = clock;
  assign uIntergerRS__reset = reset;
  assign uIntergerRS__io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uIntergerRS__io_enq = decoder_if_inst_valid & _GEN_2419; 
  assign uIntergerRS__io_enq_data = {uIntergerRS_io_enq_data_hi,uIntergerRS_io_enq_data_lo}; 
  assign uIntergerRS__io_deq = |uIntergerRS__io_deq_cond; 
  assign uIntergerRS__io_deq_cond = {uIntergerRS_io_deq_cond_hi,uIntergerRS_io_deq_cond_lo}; 
  assign uIntergerRS__io_update_entry = {uIntergerRS_io_update_entry_hi,uIntergerRS_io_update_entry_lo}; 
  assign uIntergerRS__io_update_entry_data = {uIntergerRS_io_update_entry_data_hi,uIntergerRS_io_update_entry_data_lo}; 
  assign uMulDivRS__clock = clock;
  assign uMulDivRS__reset = reset;
  assign uMulDivRS__io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uMulDivRS__io_enq = decoder_if_inst_valid & _GEN_2498; 
  assign uMulDivRS__io_enq_data = {uMulDivRS_io_enq_data_hi,uMulDivRS_io_enq_data_lo}; 
  assign uMulDivRS__io_deq = uMulDivOp_io_in_valid; 
  assign uMulDivRS__io_update_entry = {uMulDivRS_io_update_entry_hi,uMulDivRS_io_update_entry_lo}; 
  assign uMulDivRS__io_update_entry_data = {uMulDivRS_io_update_entry_data_hi,uMulDivRS_io_update_entry_data_lo}; 
  assign uLoadStoreRS__clock = clock;
  assign uLoadStoreRS__reset = reset;
  assign uLoadStoreRS__io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uLoadStoreRS__io_enq = decoder_if_inst_valid & _GEN_2490; 
  assign uLoadStoreRS__io_enq_data = {uLoadStoreRS_io_enq_data_hi,uLoadStoreRS_io_enq_data_lo}; 
  assign uLoadStoreRS__io_deq = datamem_if_ld_valid | set_ROB_store_ready; 
  assign uLoadStoreRS__io_update_entry = {uLoadStoreRS_io_update_entry_hi,uLoadStoreRS_io_update_entry_lo}; 
  assign uLoadStoreRS__io_update_entry_data = {uLoadStoreRS_io_update_entry_data_hi,uLoadStoreRS_io_update_entry_data_lo
    }; 
  assign uROB__clock = clock;
  assign uROB__reset = reset;
  assign uROB__io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uROB__io_enq = decoder_if_inst_valid & _GEN_2415; 
  assign uROB__io_enq_data = {uROB_io_enq_data_hi,33'h0}; 
  assign uROB__io_deq = uROB_io_deq_data_rob_ready & ~uROB__io_empty; 
  assign uROB__io_update_entry = {uROB_io_update_entry_hi,uROB_io_update_entry_lo}; 
  assign uROB__io_update_entry_data = {uROB_io_update_entry_data_hi,uROB_io_update_entry_data_lo}; 
  assign uCDB_clock = clock;
  assign uCDB_reset = reset;
  assign uCDB_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uCDB_io_int_valid = uIntOp_io_out_valid; 
  assign uCDB_io_int_result = uIntOp_io_out_result; 
  assign uCDB_io_int_dest = uIntOp_io_out_dest; 
  assign uCDB_io_muldiv_valid = uMulDivOp_io_out_valid; 
  assign uCDB_io_muldiv_result = uMulDivOp_io_out_result; 
  assign uCDB_io_muldiv_dest = uMulDivOp_io_out_dest; 
  assign uCDB_io_mem_valid = datamem_if_ld_data_valid; 
  assign uCDB_io_mem_result = datamem_if_ld_data; 
  assign uCDB_io_mem_dest = datamem_if_RS_idx_o; 
  assign uIntOp_clock = clock;
  assign uIntOp_reset = reset;
  assign uIntOp_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uIntOp_io_in_valid = uIntergerRS__io_deq; 
  assign uIntOp_io_in_in1 = uIntergerRS__io_deq_data[64:33]; 
  assign uIntOp_io_in_in2 = uIntergerRS__io_deq_data[32:1]; 
  assign uIntOp_io_in_op_store = uIntergerRS_io_deq_data_op[19]; 
  assign uIntOp_io_in_op_load = uIntergerRS_io_deq_data_op[18]; 
  assign uIntOp_io_in_op_muldivb_s = uIntergerRS_io_deq_data_op[17]; 
  assign uIntOp_io_in_op_muldiva_s = uIntergerRS_io_deq_data_op[16]; 
  assign uIntOp_io_in_op_div = uIntergerRS_io_deq_data_op[15]; 
  assign uIntOp_io_in_op_mul = uIntergerRS_io_deq_data_op[14]; 
  assign uIntOp_io_in_op_equal = uIntergerRS_io_deq_data_op[13]; 
  assign uIntOp_io_in_op_large = uIntergerRS_io_deq_data_op[12]; 
  assign uIntOp_io_in_op_less = uIntergerRS_io_deq_data_op[11]; 
  assign uIntOp_io_in_op_jr = uIntergerRS_io_deq_data_op[10]; 
  assign uIntOp_io_in_op_br = uIntergerRS_io_deq_data_op[9]; 
  assign uIntOp_io_in_op_sra = uIntergerRS_io_deq_data_op[8]; 
  assign uIntOp_io_in_op_srl = uIntergerRS_io_deq_data_op[7]; 
  assign uIntOp_io_in_op_sll = uIntergerRS_io_deq_data_op[6]; 
  assign uIntOp_io_in_op_sub = uIntergerRS_io_deq_data_op[5]; 
  assign uIntOp_io_in_op_add = uIntergerRS_io_deq_data_op[4]; 
  assign uIntOp_io_in_op_set = uIntergerRS_io_deq_data_op[3]; 
  assign uIntOp_io_in_op_xor = uIntergerRS_io_deq_data_op[2]; 
  assign uIntOp_io_in_op_or = uIntergerRS_io_deq_data_op[1]; 
  assign uIntOp_io_in_op_and = uIntergerRS_io_deq_data_op[0]; 
  assign uIntOp_io_in_dest = uIntergerRS__io_deq_data[111:107]; 
  assign uMulDivOp_clock = clock;
  assign uMulDivOp_reset = reset;
  assign uMulDivOp_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uMulDivOp_io_in_valid = _uMulDivOp_io_in_valid_T_4 & _uMulDivOp_io_in_valid_T_6; 
  assign uMulDivOp_io_in_in1 = uMulDivRS__io_deq_data[64:33]; 
  assign uMulDivOp_io_in_in2 = uMulDivRS__io_deq_data[32:1]; 
  assign uMulDivOp_io_in_op_muldivb_s = uMulDivRS_io_deq_data_op[17]; 
  assign uMulDivOp_io_in_op_muldiva_s = uMulDivRS_io_deq_data_op[16]; 
  assign uMulDivOp_io_in_op_mul = uMulDivRS_io_deq_data_op[14]; 
  assign uMulDivOp_io_in_dest = uMulDivRS__io_deq_data[111:107]; 
  assign uRegFile_0_clock = clock;
  assign uRegFile_0_reset = reset;
  assign uRegFile_0_io_d = 32'h0; 
  assign uRegFile_0_io_clear = 1'h1; 
  assign uRegFile_1_clock = clock;
  assign uRegFile_1_reset = reset;
  assign uRegFile_1_io_d = _T_644 ? uROB_io_deq_data_rob_value : uRegFile_io_1_q; 
  assign uRegFile_1_io_clear = 1'h0; 
  assign uRegFile_2_clock = clock;
  assign uRegFile_2_reset = reset;
  assign uRegFile_2_io_d = _T_651 ? uROB_io_deq_data_rob_value : uRegFile_io_2_q; 
  assign uRegFile_2_io_clear = 1'h0; 
  assign uRegFile_3_clock = clock;
  assign uRegFile_3_reset = reset;
  assign uRegFile_3_io_d = _T_658 ? uROB_io_deq_data_rob_value : uRegFile_io_3_q; 
  assign uRegFile_3_io_clear = 1'h0; 
  assign uRegFile_4_clock = clock;
  assign uRegFile_4_reset = reset;
  assign uRegFile_4_io_d = _T_665 ? uROB_io_deq_data_rob_value : uRegFile_io_4_q; 
  assign uRegFile_4_io_clear = 1'h0; 
  assign uRegFile_5_clock = clock;
  assign uRegFile_5_reset = reset;
  assign uRegFile_5_io_d = _T_672 ? uROB_io_deq_data_rob_value : uRegFile_io_5_q; 
  assign uRegFile_5_io_clear = 1'h0; 
  assign uRegFile_6_clock = clock;
  assign uRegFile_6_reset = reset;
  assign uRegFile_6_io_d = _T_679 ? uROB_io_deq_data_rob_value : uRegFile_io_6_q; 
  assign uRegFile_6_io_clear = 1'h0; 
  assign uRegFile_7_clock = clock;
  assign uRegFile_7_reset = reset;
  assign uRegFile_7_io_d = _T_686 ? uROB_io_deq_data_rob_value : uRegFile_io_7_q; 
  assign uRegFile_7_io_clear = 1'h0; 
  assign uRegFile_8_clock = clock;
  assign uRegFile_8_reset = reset;
  assign uRegFile_8_io_d = _T_693 ? uROB_io_deq_data_rob_value : uRegFile_io_8_q; 
  assign uRegFile_8_io_clear = 1'h0; 
  assign uRegFile_9_clock = clock;
  assign uRegFile_9_reset = reset;
  assign uRegFile_9_io_d = _T_700 ? uROB_io_deq_data_rob_value : uRegFile_io_9_q; 
  assign uRegFile_9_io_clear = 1'h0; 
  assign uRegFile_10_clock = clock;
  assign uRegFile_10_reset = reset;
  assign uRegFile_10_io_d = _T_707 ? uROB_io_deq_data_rob_value : uRegFile_io_10_q; 
  assign uRegFile_10_io_clear = 1'h0; 
  assign uRegFile_11_clock = clock;
  assign uRegFile_11_reset = reset;
  assign uRegFile_11_io_d = _T_714 ? uROB_io_deq_data_rob_value : uRegFile_io_11_q; 
  assign uRegFile_11_io_clear = 1'h0; 
  assign uRegFile_12_clock = clock;
  assign uRegFile_12_reset = reset;
  assign uRegFile_12_io_d = _T_721 ? uROB_io_deq_data_rob_value : uRegFile_io_12_q; 
  assign uRegFile_12_io_clear = 1'h0; 
  assign uRegFile_13_clock = clock;
  assign uRegFile_13_reset = reset;
  assign uRegFile_13_io_d = _T_728 ? uROB_io_deq_data_rob_value : uRegFile_io_13_q; 
  assign uRegFile_13_io_clear = 1'h0; 
  assign uRegFile_14_clock = clock;
  assign uRegFile_14_reset = reset;
  assign uRegFile_14_io_d = _T_735 ? uROB_io_deq_data_rob_value : uRegFile_io_14_q; 
  assign uRegFile_14_io_clear = 1'h0; 
  assign uRegFile_15_clock = clock;
  assign uRegFile_15_reset = reset;
  assign uRegFile_15_io_d = _T_742 ? uROB_io_deq_data_rob_value : uRegFile_io_15_q; 
  assign uRegFile_15_io_clear = 1'h0; 
  assign uRegFile_16_clock = clock;
  assign uRegFile_16_reset = reset;
  assign uRegFile_16_io_d = _T_749 ? uROB_io_deq_data_rob_value : uRegFile_io_16_q; 
  assign uRegFile_16_io_clear = 1'h0; 
  assign uRegFile_17_clock = clock;
  assign uRegFile_17_reset = reset;
  assign uRegFile_17_io_d = _T_756 ? uROB_io_deq_data_rob_value : uRegFile_io_17_q; 
  assign uRegFile_17_io_clear = 1'h0; 
  assign uRegFile_18_clock = clock;
  assign uRegFile_18_reset = reset;
  assign uRegFile_18_io_d = _T_763 ? uROB_io_deq_data_rob_value : uRegFile_io_18_q; 
  assign uRegFile_18_io_clear = 1'h0; 
  assign uRegFile_19_clock = clock;
  assign uRegFile_19_reset = reset;
  assign uRegFile_19_io_d = _T_770 ? uROB_io_deq_data_rob_value : uRegFile_io_19_q; 
  assign uRegFile_19_io_clear = 1'h0; 
  assign uRegFile_20_clock = clock;
  assign uRegFile_20_reset = reset;
  assign uRegFile_20_io_d = _T_777 ? uROB_io_deq_data_rob_value : uRegFile_io_20_q; 
  assign uRegFile_20_io_clear = 1'h0; 
  assign uRegFile_21_clock = clock;
  assign uRegFile_21_reset = reset;
  assign uRegFile_21_io_d = _T_784 ? uROB_io_deq_data_rob_value : uRegFile_io_21_q; 
  assign uRegFile_21_io_clear = 1'h0; 
  assign uRegFile_22_clock = clock;
  assign uRegFile_22_reset = reset;
  assign uRegFile_22_io_d = _T_791 ? uROB_io_deq_data_rob_value : uRegFile_io_22_q; 
  assign uRegFile_22_io_clear = 1'h0; 
  assign uRegFile_23_clock = clock;
  assign uRegFile_23_reset = reset;
  assign uRegFile_23_io_d = _T_798 ? uROB_io_deq_data_rob_value : uRegFile_io_23_q; 
  assign uRegFile_23_io_clear = 1'h0; 
  assign uRegFile_24_clock = clock;
  assign uRegFile_24_reset = reset;
  assign uRegFile_24_io_d = _T_805 ? uROB_io_deq_data_rob_value : uRegFile_io_24_q; 
  assign uRegFile_24_io_clear = 1'h0; 
  assign uRegFile_25_clock = clock;
  assign uRegFile_25_reset = reset;
  assign uRegFile_25_io_d = _T_812 ? uROB_io_deq_data_rob_value : uRegFile_io_25_q; 
  assign uRegFile_25_io_clear = 1'h0; 
  assign uRegFile_26_clock = clock;
  assign uRegFile_26_reset = reset;
  assign uRegFile_26_io_d = _T_819 ? uROB_io_deq_data_rob_value : uRegFile_io_26_q; 
  assign uRegFile_26_io_clear = 1'h0; 
  assign uRegFile_27_clock = clock;
  assign uRegFile_27_reset = reset;
  assign uRegFile_27_io_d = _T_826 ? uROB_io_deq_data_rob_value : uRegFile_io_27_q; 
  assign uRegFile_27_io_clear = 1'h0; 
  assign uRegFile_28_clock = clock;
  assign uRegFile_28_reset = reset;
  assign uRegFile_28_io_d = _T_833 ? uROB_io_deq_data_rob_value : uRegFile_io_28_q; 
  assign uRegFile_28_io_clear = 1'h0; 
  assign uRegFile_29_clock = clock;
  assign uRegFile_29_reset = reset;
  assign uRegFile_29_io_d = _T_840 ? uROB_io_deq_data_rob_value : uRegFile_io_29_q; 
  assign uRegFile_29_io_clear = 1'h0; 
  assign uRegFile_30_clock = clock;
  assign uRegFile_30_reset = reset;
  assign uRegFile_30_io_d = _T_847 ? uROB_io_deq_data_rob_value : uRegFile_io_30_q; 
  assign uRegFile_30_io_clear = 1'h0; 
  assign uRegFile_31_clock = clock;
  assign uRegFile_31_reset = reset;
  assign uRegFile_31_io_d = _T_854 ? uROB_io_deq_data_rob_value : uRegFile_io_31_q; 
  assign uRegFile_31_io_clear = 1'h0; 
  assign uRegState_0_clock = clock;
  assign uRegState_0_reset = reset;
  assign uRegState_0_io_d_busy = decoder_if_inst_valid ? _GEN_2458 : _GEN_21; 
  assign uRegState_0_io_d_reorder = decoder_if_inst_valid ? _GEN_2426 : _GEN_20; 
  assign uRegState_0_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_1_clock = clock;
  assign uRegState_1_reset = reset;
  assign uRegState_1_io_d_busy = decoder_if_inst_valid ? _GEN_2459 : _GEN_23; 
  assign uRegState_1_io_d_reorder = decoder_if_inst_valid ? _GEN_2427 : _GEN_22; 
  assign uRegState_1_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_2_clock = clock;
  assign uRegState_2_reset = reset;
  assign uRegState_2_io_d_busy = decoder_if_inst_valid ? _GEN_2460 : _GEN_25; 
  assign uRegState_2_io_d_reorder = decoder_if_inst_valid ? _GEN_2428 : _GEN_24; 
  assign uRegState_2_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_3_clock = clock;
  assign uRegState_3_reset = reset;
  assign uRegState_3_io_d_busy = decoder_if_inst_valid ? _GEN_2461 : _GEN_27; 
  assign uRegState_3_io_d_reorder = decoder_if_inst_valid ? _GEN_2429 : _GEN_26; 
  assign uRegState_3_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_4_clock = clock;
  assign uRegState_4_reset = reset;
  assign uRegState_4_io_d_busy = decoder_if_inst_valid ? _GEN_2462 : _GEN_29; 
  assign uRegState_4_io_d_reorder = decoder_if_inst_valid ? _GEN_2430 : _GEN_28; 
  assign uRegState_4_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_5_clock = clock;
  assign uRegState_5_reset = reset;
  assign uRegState_5_io_d_busy = decoder_if_inst_valid ? _GEN_2463 : _GEN_31; 
  assign uRegState_5_io_d_reorder = decoder_if_inst_valid ? _GEN_2431 : _GEN_30; 
  assign uRegState_5_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_6_clock = clock;
  assign uRegState_6_reset = reset;
  assign uRegState_6_io_d_busy = decoder_if_inst_valid ? _GEN_2464 : _GEN_33; 
  assign uRegState_6_io_d_reorder = decoder_if_inst_valid ? _GEN_2432 : _GEN_32; 
  assign uRegState_6_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_7_clock = clock;
  assign uRegState_7_reset = reset;
  assign uRegState_7_io_d_busy = decoder_if_inst_valid ? _GEN_2465 : _GEN_35; 
  assign uRegState_7_io_d_reorder = decoder_if_inst_valid ? _GEN_2433 : _GEN_34; 
  assign uRegState_7_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_8_clock = clock;
  assign uRegState_8_reset = reset;
  assign uRegState_8_io_d_busy = decoder_if_inst_valid ? _GEN_2466 : _GEN_37; 
  assign uRegState_8_io_d_reorder = decoder_if_inst_valid ? _GEN_2434 : _GEN_36; 
  assign uRegState_8_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_9_clock = clock;
  assign uRegState_9_reset = reset;
  assign uRegState_9_io_d_busy = decoder_if_inst_valid ? _GEN_2467 : _GEN_39; 
  assign uRegState_9_io_d_reorder = decoder_if_inst_valid ? _GEN_2435 : _GEN_38; 
  assign uRegState_9_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_10_clock = clock;
  assign uRegState_10_reset = reset;
  assign uRegState_10_io_d_busy = decoder_if_inst_valid ? _GEN_2468 : _GEN_41; 
  assign uRegState_10_io_d_reorder = decoder_if_inst_valid ? _GEN_2436 : _GEN_40; 
  assign uRegState_10_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_11_clock = clock;
  assign uRegState_11_reset = reset;
  assign uRegState_11_io_d_busy = decoder_if_inst_valid ? _GEN_2469 : _GEN_43; 
  assign uRegState_11_io_d_reorder = decoder_if_inst_valid ? _GEN_2437 : _GEN_42; 
  assign uRegState_11_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_12_clock = clock;
  assign uRegState_12_reset = reset;
  assign uRegState_12_io_d_busy = decoder_if_inst_valid ? _GEN_2470 : _GEN_45; 
  assign uRegState_12_io_d_reorder = decoder_if_inst_valid ? _GEN_2438 : _GEN_44; 
  assign uRegState_12_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_13_clock = clock;
  assign uRegState_13_reset = reset;
  assign uRegState_13_io_d_busy = decoder_if_inst_valid ? _GEN_2471 : _GEN_47; 
  assign uRegState_13_io_d_reorder = decoder_if_inst_valid ? _GEN_2439 : _GEN_46; 
  assign uRegState_13_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_14_clock = clock;
  assign uRegState_14_reset = reset;
  assign uRegState_14_io_d_busy = decoder_if_inst_valid ? _GEN_2472 : _GEN_49; 
  assign uRegState_14_io_d_reorder = decoder_if_inst_valid ? _GEN_2440 : _GEN_48; 
  assign uRegState_14_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_15_clock = clock;
  assign uRegState_15_reset = reset;
  assign uRegState_15_io_d_busy = decoder_if_inst_valid ? _GEN_2473 : _GEN_51; 
  assign uRegState_15_io_d_reorder = decoder_if_inst_valid ? _GEN_2441 : _GEN_50; 
  assign uRegState_15_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_16_clock = clock;
  assign uRegState_16_reset = reset;
  assign uRegState_16_io_d_busy = decoder_if_inst_valid ? _GEN_2474 : _GEN_53; 
  assign uRegState_16_io_d_reorder = decoder_if_inst_valid ? _GEN_2442 : _GEN_52; 
  assign uRegState_16_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_17_clock = clock;
  assign uRegState_17_reset = reset;
  assign uRegState_17_io_d_busy = decoder_if_inst_valid ? _GEN_2475 : _GEN_55; 
  assign uRegState_17_io_d_reorder = decoder_if_inst_valid ? _GEN_2443 : _GEN_54; 
  assign uRegState_17_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_18_clock = clock;
  assign uRegState_18_reset = reset;
  assign uRegState_18_io_d_busy = decoder_if_inst_valid ? _GEN_2476 : _GEN_57; 
  assign uRegState_18_io_d_reorder = decoder_if_inst_valid ? _GEN_2444 : _GEN_56; 
  assign uRegState_18_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_19_clock = clock;
  assign uRegState_19_reset = reset;
  assign uRegState_19_io_d_busy = decoder_if_inst_valid ? _GEN_2477 : _GEN_59; 
  assign uRegState_19_io_d_reorder = decoder_if_inst_valid ? _GEN_2445 : _GEN_58; 
  assign uRegState_19_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_20_clock = clock;
  assign uRegState_20_reset = reset;
  assign uRegState_20_io_d_busy = decoder_if_inst_valid ? _GEN_2478 : _GEN_61; 
  assign uRegState_20_io_d_reorder = decoder_if_inst_valid ? _GEN_2446 : _GEN_60; 
  assign uRegState_20_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_21_clock = clock;
  assign uRegState_21_reset = reset;
  assign uRegState_21_io_d_busy = decoder_if_inst_valid ? _GEN_2479 : _GEN_63; 
  assign uRegState_21_io_d_reorder = decoder_if_inst_valid ? _GEN_2447 : _GEN_62; 
  assign uRegState_21_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_22_clock = clock;
  assign uRegState_22_reset = reset;
  assign uRegState_22_io_d_busy = decoder_if_inst_valid ? _GEN_2480 : _GEN_65; 
  assign uRegState_22_io_d_reorder = decoder_if_inst_valid ? _GEN_2448 : _GEN_64; 
  assign uRegState_22_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_23_clock = clock;
  assign uRegState_23_reset = reset;
  assign uRegState_23_io_d_busy = decoder_if_inst_valid ? _GEN_2481 : _GEN_67; 
  assign uRegState_23_io_d_reorder = decoder_if_inst_valid ? _GEN_2449 : _GEN_66; 
  assign uRegState_23_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_24_clock = clock;
  assign uRegState_24_reset = reset;
  assign uRegState_24_io_d_busy = decoder_if_inst_valid ? _GEN_2482 : _GEN_69; 
  assign uRegState_24_io_d_reorder = decoder_if_inst_valid ? _GEN_2450 : _GEN_68; 
  assign uRegState_24_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_25_clock = clock;
  assign uRegState_25_reset = reset;
  assign uRegState_25_io_d_busy = decoder_if_inst_valid ? _GEN_2483 : _GEN_71; 
  assign uRegState_25_io_d_reorder = decoder_if_inst_valid ? _GEN_2451 : _GEN_70; 
  assign uRegState_25_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_26_clock = clock;
  assign uRegState_26_reset = reset;
  assign uRegState_26_io_d_busy = decoder_if_inst_valid ? _GEN_2484 : _GEN_73; 
  assign uRegState_26_io_d_reorder = decoder_if_inst_valid ? _GEN_2452 : _GEN_72; 
  assign uRegState_26_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_27_clock = clock;
  assign uRegState_27_reset = reset;
  assign uRegState_27_io_d_busy = decoder_if_inst_valid ? _GEN_2485 : _GEN_75; 
  assign uRegState_27_io_d_reorder = decoder_if_inst_valid ? _GEN_2453 : _GEN_74; 
  assign uRegState_27_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_28_clock = clock;
  assign uRegState_28_reset = reset;
  assign uRegState_28_io_d_busy = decoder_if_inst_valid ? _GEN_2486 : _GEN_77; 
  assign uRegState_28_io_d_reorder = decoder_if_inst_valid ? _GEN_2454 : _GEN_76; 
  assign uRegState_28_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_29_clock = clock;
  assign uRegState_29_reset = reset;
  assign uRegState_29_io_d_busy = decoder_if_inst_valid ? _GEN_2487 : _GEN_79; 
  assign uRegState_29_io_d_reorder = decoder_if_inst_valid ? _GEN_2455 : _GEN_78; 
  assign uRegState_29_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_30_clock = clock;
  assign uRegState_30_reset = reset;
  assign uRegState_30_io_d_busy = decoder_if_inst_valid ? _GEN_2488 : _GEN_81; 
  assign uRegState_30_io_d_reorder = decoder_if_inst_valid ? _GEN_2456 : _GEN_80; 
  assign uRegState_30_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uRegState_31_clock = clock;
  assign uRegState_31_reset = reset;
  assign uRegState_31_io_d_busy = decoder_if_inst_valid ? _GEN_2489 : _GEN_83; 
  assign uRegState_31_io_d_reorder = decoder_if_inst_valid ? _GEN_2457 : _GEN_82; 
  assign uRegState_31_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign integer_inst_r_clock = clock;
  assign integer_inst_r_reset = reset;
  assign integer_inst_r_io_d = _integer_inst_r_io_d_T_13 | _integer_inst_r_io_d_T_15; 
  assign integer_inst_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign branch_inst_r_clock = clock;
  assign branch_inst_r_reset = reset;
  assign branch_inst_r_io_d = decoder_if_exe_op_br; 
  assign branch_inst_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign store_inst_r_clock = clock;
  assign store_inst_r_reset = reset;
  assign store_inst_r_io_d = decoder_if_exe_op_store; 
  assign store_inst_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign load_inst_r_clock = clock;
  assign load_inst_r_reset = reset;
  assign load_inst_r_io_d = decoder_if_exe_op_load; 
  assign load_inst_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign muldiv_inst_r_clock = clock;
  assign muldiv_inst_r_reset = reset;
  assign muldiv_inst_r_io_d = decoder_if_exe_op_mul | decoder_if_exe_op_div; 
  assign muldiv_inst_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign mBranchProc_st_clock = clock;
  assign mBranchProc_st_reset = reset;
  assign mBranchProc_st_io_d = 2'h0 == branchProc_stEnum ? _GEN_13 : _GEN_17; 
  assign mBranchProc_st_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign re_jump_addr_r_clock = clock;
  assign re_jump_addr_r_reset = reset;
  assign re_jump_addr_r_io_d = uROB_io_deq_data_rob_ready ? _GEN_2978 : re_jump_addr_r_io_q; 
  assign re_jump_addr_r_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uIntBusGetData_st_clock = clock;
  assign uIntBusGetData_st_reset = reset;
  assign uIntBusGetData_st_io_d = uIntBusGetData_st_io_q ? ~uCDB_io_int_ready : uIntOp_io_in_valid; 
  assign uIntBusGetData_st_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uMulDivBusGetData_st_clock = clock;
  assign uMulDivBusGetData_st_reset = reset;
  assign uMulDivBusGetData_st_io_d = uMulDivBusGetData_st_io_q ? ~uCDB_io_muldiv_ready : uMulDivOp_io_in_valid; 
  assign uMulDivBusGetData_st_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
  assign uLoadBusGetData_st_clock = clock;
  assign uLoadBusGetData_st_reset = reset;
  assign uLoadBusGetData_st_io_d = uLoadBusGetData_st_io_q ? ~uCDB_io_mem_ready : datamem_if_ld_valid; 
  assign uLoadBusGetData_st_io_clear = uROB_io_deq_data_rob_ready & _GEN_2979; 
endmodule
